-- nios_system.vhd

-- Generated using ACDS version 13.0sp1 232 at 2019.10.18.16:55:22

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity nios_system is
	port (
		zs_addr_from_the_SDRAM      : out   std_logic_vector(12 downto 0);                    --       SDRAM_wire.addr
		zs_ba_from_the_SDRAM        : out   std_logic_vector(1 downto 0);                     --                 .ba
		zs_cas_n_from_the_SDRAM     : out   std_logic;                                        --                 .cas_n
		zs_cke_from_the_SDRAM       : out   std_logic;                                        --                 .cke
		zs_cs_n_from_the_SDRAM      : out   std_logic;                                        --                 .cs_n
		zs_dq_to_and_from_the_SDRAM : inout std_logic_vector(15 downto 0) := (others => '0'); --                 .dq
		zs_dqm_from_the_SDRAM       : out   std_logic_vector(1 downto 0);                     --                 .dqm
		zs_ras_n_from_the_SDRAM     : out   std_logic;                                        --                 .ras_n
		zs_we_n_from_the_SDRAM      : out   std_logic;                                        --                 .we_n
		reset_n                     : in    std_logic                     := '0';             -- clk_clk_in_reset.reset_n
		clk                         : in    std_logic                     := '0';             --       clk_clk_in.clk
		sdram_clk                   : out   std_logic;                                        --            sdram.clk
		omoteurctr_export           : out   std_logic_vector(31 downto 0);                    --       omoteurctr.export
		capt3_0_signal_export       : in    std_logic_vector(31 downto 0) := (others => '0'); --   capt3_0_signal.export
		capt6_4_signal_export       : in    std_logic_vector(31 downto 0) := (others => '0')  --   capt6_4_signal.export
	);
end entity nios_system;

architecture rtl of nios_system is
	component nios_system_JTAG_UART is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component nios_system_JTAG_UART;

	component nios_system_Interval_timer is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component nios_system_Interval_timer;

	component nios_system_SDRAM is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(23 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(12 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component nios_system_SDRAM;

	component nios_system_CPU is
		port (
			clk                                   : in  std_logic                     := 'X';             -- clk
			reset_n                               : in  std_logic                     := 'X';             -- reset_n
			d_address                             : out std_logic_vector(28 downto 0);                    -- address
			d_byteenable                          : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                                : out std_logic;                                        -- read
			d_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_write                               : out std_logic;                                        -- write
			d_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_debug_module_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                             : out std_logic_vector(27 downto 0);                    -- address
			i_read                                : out std_logic;                                        -- read
			i_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                       : in  std_logic                     := 'X';             -- readdatavalid
			d_irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			jtag_debug_module_resetrequest        : out std_logic;                                        -- reset
			jtag_debug_module_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			jtag_debug_module_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			jtag_debug_module_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			jtag_debug_module_read                : in  std_logic                     := 'X';             -- read
			jtag_debug_module_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			jtag_debug_module_waitrequest         : out std_logic;                                        -- waitrequest
			jtag_debug_module_write               : in  std_logic                     := 'X';             -- write
			jtag_debug_module_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			no_ci_readra                          : out std_logic                                         -- readra
		);
	end component nios_system_CPU;

	component nios_system_sysid is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component nios_system_sysid;

	component nios_system_External_Clocks is
		port (
			CLOCK_50    : in  std_logic := 'X'; -- clk
			reset       : in  std_logic := 'X'; -- reset
			sys_clk     : out std_logic;        -- clk
			sys_reset_n : out std_logic;        -- reset_n
			SDRAM_CLK   : out std_logic         -- clk
		);
	end component nios_system_External_Clocks;

	component nios_system_CTR_MOTEUR is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset      : in  std_logic                     := 'X';             -- reset
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			chipselect : in  std_logic                     := 'X';             -- chipselect
			read       : in  std_logic                     := 'X';             -- read
			write      : in  std_logic                     := 'X';             -- write
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(31 downto 0)                     -- export
		);
	end component nios_system_CTR_MOTEUR;

	component nios_system_capt3_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset      : in  std_logic                     := 'X';             -- reset
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			chipselect : in  std_logic                     := 'X';             -- chipselect
			read       : in  std_logic                     := 'X';             -- read
			write      : in  std_logic                     := 'X';             -- write
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(31 downto 0) := (others => 'X')  -- export
		);
	end component nios_system_capt3_0;

	component altera_merlin_master_agent is
		generic (
			PKT_PROTECTION_H          : integer := 80;
			PKT_PROTECTION_L          : integer := 80;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_BURSTWRAP_H           : integer := 79;
			PKT_BURSTWRAP_L           : integer := 77;
			PKT_BURST_SIZE_H          : integer := 86;
			PKT_BURST_SIZE_L          : integer := 84;
			PKT_BURST_TYPE_H          : integer := 94;
			PKT_BURST_TYPE_L          : integer := 93;
			PKT_BYTE_CNT_H            : integer := 76;
			PKT_BYTE_CNT_L            : integer := 74;
			PKT_ADDR_H                : integer := 73;
			PKT_ADDR_L                : integer := 42;
			PKT_TRANS_COMPRESSED_READ : integer := 41;
			PKT_TRANS_POSTED          : integer := 40;
			PKT_TRANS_WRITE           : integer := 39;
			PKT_TRANS_READ            : integer := 38;
			PKT_TRANS_LOCK            : integer := 82;
			PKT_TRANS_EXCLUSIVE       : integer := 83;
			PKT_DATA_H                : integer := 37;
			PKT_DATA_L                : integer := 6;
			PKT_BYTEEN_H              : integer := 5;
			PKT_BYTEEN_L              : integer := 2;
			PKT_SRC_ID_H              : integer := 1;
			PKT_SRC_ID_L              : integer := 1;
			PKT_DEST_ID_H             : integer := 0;
			PKT_DEST_ID_L             : integer := 0;
			PKT_THREAD_ID_H           : integer := 88;
			PKT_THREAD_ID_L           : integer := 87;
			PKT_CACHE_H               : integer := 92;
			PKT_CACHE_L               : integer := 89;
			PKT_DATA_SIDEBAND_H       : integer := 105;
			PKT_DATA_SIDEBAND_L       : integer := 98;
			PKT_QOS_H                 : integer := 109;
			PKT_QOS_L                 : integer := 106;
			PKT_ADDR_SIDEBAND_H       : integer := 97;
			PKT_ADDR_SIDEBAND_L       : integer := 93;
			PKT_RESPONSE_STATUS_H     : integer := 111;
			PKT_RESPONSE_STATUS_L     : integer := 110;
			ST_DATA_W                 : integer := 112;
			ST_CHANNEL_W              : integer := 1;
			AV_BURSTCOUNT_W           : integer := 3;
			SUPPRESS_0_BYTEEN_RSP     : integer := 1;
			ID                        : integer := 1;
			BURSTWRAP_VALUE           : integer := 4;
			CACHE_VALUE               : integer := 0;
			SECURE_ACCESS_BIT         : integer := 1;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                      := 'X';             -- clk
			reset                   : in  std_logic                      := 'X';             -- reset
			av_address              : in  std_logic_vector(28 downto 0)  := (others => 'X'); -- address
			av_write                : in  std_logic                      := 'X';             -- write
			av_read                 : in  std_logic                      := 'X';             -- read
			av_writedata            : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			av_readdata             : out std_logic_vector(31 downto 0);                     -- readdata
			av_waitrequest          : out std_logic;                                         -- waitrequest
			av_readdatavalid        : out std_logic;                                         -- readdatavalid
			av_byteenable           : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			av_burstcount           : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- burstcount
			av_debugaccess          : in  std_logic                      := 'X';             -- debugaccess
			av_lock                 : in  std_logic                      := 'X';             -- lock
			cp_valid                : out std_logic;                                         -- valid
			cp_data                 : out std_logic_vector(101 downto 0);                    -- data
			cp_startofpacket        : out std_logic;                                         -- startofpacket
			cp_endofpacket          : out std_logic;                                         -- endofpacket
			cp_ready                : in  std_logic                      := 'X';             -- ready
			rp_valid                : in  std_logic                      := 'X';             -- valid
			rp_data                 : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			rp_channel              : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- channel
			rp_startofpacket        : in  std_logic                      := 'X';             -- startofpacket
			rp_endofpacket          : in  std_logic                      := 'X';             -- endofpacket
			rp_ready                : out std_logic;                                         -- ready
			av_response             : out std_logic_vector(1 downto 0);                      -- response
			av_writeresponserequest : in  std_logic                      := 'X';             -- writeresponserequest
			av_writeresponsevalid   : out std_logic                                          -- writeresponsevalid
		);
	end component altera_merlin_master_agent;

	component nios_system_addr_router is
		port (
			sink_ready         : out std_logic;                                         -- ready
			sink_valid         : in  std_logic                      := 'X';             -- valid
			sink_data          : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			src_ready          : in  std_logic                      := 'X';             -- ready
			src_valid          : out std_logic;                                         -- valid
			src_data           : out std_logic_vector(101 downto 0);                    -- data
			src_channel        : out std_logic_vector(7 downto 0);                      -- channel
			src_startofpacket  : out std_logic;                                         -- startofpacket
			src_endofpacket    : out std_logic                                          -- endofpacket
		);
	end component nios_system_addr_router;

	component nios_system_addr_router_001 is
		port (
			sink_ready         : out std_logic;                                         -- ready
			sink_valid         : in  std_logic                      := 'X';             -- valid
			sink_data          : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			src_ready          : in  std_logic                      := 'X';             -- ready
			src_valid          : out std_logic;                                         -- valid
			src_data           : out std_logic_vector(101 downto 0);                    -- data
			src_channel        : out std_logic_vector(7 downto 0);                      -- channel
			src_startofpacket  : out std_logic;                                         -- startofpacket
			src_endofpacket    : out std_logic                                          -- endofpacket
		);
	end component nios_system_addr_router_001;

	component nios_system_id_router is
		port (
			sink_ready         : out std_logic;                                         -- ready
			sink_valid         : in  std_logic                      := 'X';             -- valid
			sink_data          : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			src_ready          : in  std_logic                      := 'X';             -- ready
			src_valid          : out std_logic;                                         -- valid
			src_data           : out std_logic_vector(101 downto 0);                    -- data
			src_channel        : out std_logic_vector(7 downto 0);                      -- channel
			src_startofpacket  : out std_logic;                                         -- startofpacket
			src_endofpacket    : out std_logic                                          -- endofpacket
		);
	end component nios_system_id_router;

	component nios_system_id_router_001 is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(83 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(83 downto 0);                    -- data
			src_channel        : out std_logic_vector(7 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component nios_system_id_router_001;

	component nios_system_id_router_002 is
		port (
			sink_ready         : out std_logic;                                         -- ready
			sink_valid         : in  std_logic                      := 'X';             -- valid
			sink_data          : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			src_ready          : in  std_logic                      := 'X';             -- ready
			src_valid          : out std_logic;                                         -- valid
			src_data           : out std_logic_vector(101 downto 0);                    -- data
			src_channel        : out std_logic_vector(7 downto 0);                      -- channel
			src_startofpacket  : out std_logic;                                         -- startofpacket
			src_endofpacket    : out std_logic                                          -- endofpacket
		);
	end component nios_system_id_router_002;

	component altera_merlin_traffic_limiter is
		generic (
			PKT_DEST_ID_H             : integer := 0;
			PKT_DEST_ID_L             : integer := 0;
			PKT_TRANS_POSTED          : integer := 0;
			PKT_TRANS_WRITE           : integer := 0;
			MAX_OUTSTANDING_RESPONSES : integer := 0;
			PIPELINED                 : integer := 0;
			ST_DATA_W                 : integer := 72;
			ST_CHANNEL_W              : integer := 1;
			VALID_WIDTH               : integer := 1;
			ENFORCE_ORDER             : integer := 1;
			PREVENT_HAZARDS           : integer := 0;
			PKT_BYTE_CNT_H            : integer := 0;
			PKT_BYTE_CNT_L            : integer := 0;
			PKT_BYTEEN_H              : integer := 0;
			PKT_BYTEEN_L              : integer := 0
		);
		port (
			clk                    : in  std_logic                      := 'X';             -- clk
			reset                  : in  std_logic                      := 'X';             -- reset
			cmd_sink_ready         : out std_logic;                                         -- ready
			cmd_sink_valid         : in  std_logic                      := 'X';             -- valid
			cmd_sink_data          : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			cmd_sink_channel       : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- channel
			cmd_sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			cmd_sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			cmd_src_ready          : in  std_logic                      := 'X';             -- ready
			cmd_src_data           : out std_logic_vector(101 downto 0);                    -- data
			cmd_src_channel        : out std_logic_vector(7 downto 0);                      -- channel
			cmd_src_startofpacket  : out std_logic;                                         -- startofpacket
			cmd_src_endofpacket    : out std_logic;                                         -- endofpacket
			rsp_sink_ready         : out std_logic;                                         -- ready
			rsp_sink_valid         : in  std_logic                      := 'X';             -- valid
			rsp_sink_channel       : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- channel
			rsp_sink_data          : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			rsp_sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			rsp_sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			rsp_src_ready          : in  std_logic                      := 'X';             -- ready
			rsp_src_valid          : out std_logic;                                         -- valid
			rsp_src_data           : out std_logic_vector(101 downto 0);                    -- data
			rsp_src_channel        : out std_logic_vector(7 downto 0);                      -- channel
			rsp_src_startofpacket  : out std_logic;                                         -- startofpacket
			rsp_src_endofpacket    : out std_logic;                                         -- endofpacket
			cmd_src_valid          : out std_logic_vector(7 downto 0)                       -- data
		);
	end component altera_merlin_traffic_limiter;

	component altera_merlin_burst_adapter is
		generic (
			PKT_ADDR_H                : integer := 79;
			PKT_ADDR_L                : integer := 48;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_BYTE_CNT_H            : integer := 5;
			PKT_BYTE_CNT_L            : integer := 0;
			PKT_BYTEEN_H              : integer := 83;
			PKT_BYTEEN_L              : integer := 80;
			PKT_BURST_SIZE_H          : integer := 86;
			PKT_BURST_SIZE_L          : integer := 84;
			PKT_BURST_TYPE_H          : integer := 88;
			PKT_BURST_TYPE_L          : integer := 87;
			PKT_BURSTWRAP_H           : integer := 11;
			PKT_BURSTWRAP_L           : integer := 6;
			PKT_TRANS_COMPRESSED_READ : integer := 14;
			PKT_TRANS_WRITE           : integer := 13;
			PKT_TRANS_READ            : integer := 12;
			OUT_NARROW_SIZE           : integer := 0;
			IN_NARROW_SIZE            : integer := 0;
			OUT_FIXED                 : integer := 0;
			OUT_COMPLETE_WRAP         : integer := 0;
			ST_DATA_W                 : integer := 89;
			ST_CHANNEL_W              : integer := 8;
			OUT_BYTE_CNT_H            : integer := 5;
			OUT_BURSTWRAP_H           : integer := 11;
			COMPRESSED_READ_SUPPORT   : integer := 1;
			BYTEENABLE_SYNTHESIS      : integer := 0;
			PIPE_INPUTS               : integer := 0;
			NO_WRAP_SUPPORT           : integer := 0;
			BURSTWRAP_CONST_MASK      : integer := 0;
			BURSTWRAP_CONST_VALUE     : integer := -1
		);
		port (
			clk                   : in  std_logic                     := 'X';             -- clk
			reset                 : in  std_logic                     := 'X';             -- reset
			sink0_valid           : in  std_logic                     := 'X';             -- valid
			sink0_data            : in  std_logic_vector(83 downto 0) := (others => 'X'); -- data
			sink0_channel         : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- channel
			sink0_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			sink0_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			sink0_ready           : out std_logic;                                        -- ready
			source0_valid         : out std_logic;                                        -- valid
			source0_data          : out std_logic_vector(83 downto 0);                    -- data
			source0_channel       : out std_logic_vector(7 downto 0);                     -- channel
			source0_startofpacket : out std_logic;                                        -- startofpacket
			source0_endofpacket   : out std_logic;                                        -- endofpacket
			source0_ready         : in  std_logic                     := 'X'              -- ready
		);
	end component altera_merlin_burst_adapter;

	component nios_system_cmd_xbar_demux is
		port (
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			sink_ready         : out std_logic;                                         -- ready
			sink_channel       : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- data
			src0_ready         : in  std_logic                      := 'X';             -- ready
			src0_valid         : out std_logic;                                         -- valid
			src0_data          : out std_logic_vector(101 downto 0);                    -- data
			src0_channel       : out std_logic_vector(7 downto 0);                      -- channel
			src0_startofpacket : out std_logic;                                         -- startofpacket
			src0_endofpacket   : out std_logic;                                         -- endofpacket
			src1_ready         : in  std_logic                      := 'X';             -- ready
			src1_valid         : out std_logic;                                         -- valid
			src1_data          : out std_logic_vector(101 downto 0);                    -- data
			src1_channel       : out std_logic_vector(7 downto 0);                      -- channel
			src1_startofpacket : out std_logic;                                         -- startofpacket
			src1_endofpacket   : out std_logic                                          -- endofpacket
		);
	end component nios_system_cmd_xbar_demux;

	component nios_system_cmd_xbar_demux_001 is
		port (
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			sink_ready         : out std_logic;                                         -- ready
			sink_channel       : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- valid
			src0_ready         : in  std_logic                      := 'X';             -- ready
			src0_valid         : out std_logic;                                         -- valid
			src0_data          : out std_logic_vector(101 downto 0);                    -- data
			src0_channel       : out std_logic_vector(7 downto 0);                      -- channel
			src0_startofpacket : out std_logic;                                         -- startofpacket
			src0_endofpacket   : out std_logic;                                         -- endofpacket
			src1_ready         : in  std_logic                      := 'X';             -- ready
			src1_valid         : out std_logic;                                         -- valid
			src1_data          : out std_logic_vector(101 downto 0);                    -- data
			src1_channel       : out std_logic_vector(7 downto 0);                      -- channel
			src1_startofpacket : out std_logic;                                         -- startofpacket
			src1_endofpacket   : out std_logic;                                         -- endofpacket
			src2_ready         : in  std_logic                      := 'X';             -- ready
			src2_valid         : out std_logic;                                         -- valid
			src2_data          : out std_logic_vector(101 downto 0);                    -- data
			src2_channel       : out std_logic_vector(7 downto 0);                      -- channel
			src2_startofpacket : out std_logic;                                         -- startofpacket
			src2_endofpacket   : out std_logic;                                         -- endofpacket
			src3_ready         : in  std_logic                      := 'X';             -- ready
			src3_valid         : out std_logic;                                         -- valid
			src3_data          : out std_logic_vector(101 downto 0);                    -- data
			src3_channel       : out std_logic_vector(7 downto 0);                      -- channel
			src3_startofpacket : out std_logic;                                         -- startofpacket
			src3_endofpacket   : out std_logic;                                         -- endofpacket
			src4_ready         : in  std_logic                      := 'X';             -- ready
			src4_valid         : out std_logic;                                         -- valid
			src4_data          : out std_logic_vector(101 downto 0);                    -- data
			src4_channel       : out std_logic_vector(7 downto 0);                      -- channel
			src4_startofpacket : out std_logic;                                         -- startofpacket
			src4_endofpacket   : out std_logic;                                         -- endofpacket
			src5_ready         : in  std_logic                      := 'X';             -- ready
			src5_valid         : out std_logic;                                         -- valid
			src5_data          : out std_logic_vector(101 downto 0);                    -- data
			src5_channel       : out std_logic_vector(7 downto 0);                      -- channel
			src5_startofpacket : out std_logic;                                         -- startofpacket
			src5_endofpacket   : out std_logic;                                         -- endofpacket
			src6_ready         : in  std_logic                      := 'X';             -- ready
			src6_valid         : out std_logic;                                         -- valid
			src6_data          : out std_logic_vector(101 downto 0);                    -- data
			src6_channel       : out std_logic_vector(7 downto 0);                      -- channel
			src6_startofpacket : out std_logic;                                         -- startofpacket
			src6_endofpacket   : out std_logic;                                         -- endofpacket
			src7_ready         : in  std_logic                      := 'X';             -- ready
			src7_valid         : out std_logic;                                         -- valid
			src7_data          : out std_logic_vector(101 downto 0);                    -- data
			src7_channel       : out std_logic_vector(7 downto 0);                      -- channel
			src7_startofpacket : out std_logic;                                         -- startofpacket
			src7_endofpacket   : out std_logic                                          -- endofpacket
		);
	end component nios_system_cmd_xbar_demux_001;

	component nios_system_cmd_xbar_mux is
		port (
			clk                 : in  std_logic                      := 'X';             -- clk
			reset               : in  std_logic                      := 'X';             -- reset
			src_ready           : in  std_logic                      := 'X';             -- ready
			src_valid           : out std_logic;                                         -- valid
			src_data            : out std_logic_vector(101 downto 0);                    -- data
			src_channel         : out std_logic_vector(7 downto 0);                      -- channel
			src_startofpacket   : out std_logic;                                         -- startofpacket
			src_endofpacket     : out std_logic;                                         -- endofpacket
			sink0_ready         : out std_logic;                                         -- ready
			sink0_valid         : in  std_logic                      := 'X';             -- valid
			sink0_channel       : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- channel
			sink0_data          : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink0_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink0_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink1_ready         : out std_logic;                                         -- ready
			sink1_valid         : in  std_logic                      := 'X';             -- valid
			sink1_channel       : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- channel
			sink1_data          : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink1_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink1_endofpacket   : in  std_logic                      := 'X'              -- endofpacket
		);
	end component nios_system_cmd_xbar_mux;

	component nios_system_rsp_xbar_demux is
		port (
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			sink_ready         : out std_logic;                                         -- ready
			sink_channel       : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- valid
			src0_ready         : in  std_logic                      := 'X';             -- ready
			src0_valid         : out std_logic;                                         -- valid
			src0_data          : out std_logic_vector(101 downto 0);                    -- data
			src0_channel       : out std_logic_vector(7 downto 0);                      -- channel
			src0_startofpacket : out std_logic;                                         -- startofpacket
			src0_endofpacket   : out std_logic;                                         -- endofpacket
			src1_ready         : in  std_logic                      := 'X';             -- ready
			src1_valid         : out std_logic;                                         -- valid
			src1_data          : out std_logic_vector(101 downto 0);                    -- data
			src1_channel       : out std_logic_vector(7 downto 0);                      -- channel
			src1_startofpacket : out std_logic;                                         -- startofpacket
			src1_endofpacket   : out std_logic                                          -- endofpacket
		);
	end component nios_system_rsp_xbar_demux;

	component nios_system_rsp_xbar_demux_002 is
		port (
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			sink_ready         : out std_logic;                                         -- ready
			sink_channel       : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- valid
			src0_ready         : in  std_logic                      := 'X';             -- ready
			src0_valid         : out std_logic;                                         -- valid
			src0_data          : out std_logic_vector(101 downto 0);                    -- data
			src0_channel       : out std_logic_vector(7 downto 0);                      -- channel
			src0_startofpacket : out std_logic;                                         -- startofpacket
			src0_endofpacket   : out std_logic                                          -- endofpacket
		);
	end component nios_system_rsp_xbar_demux_002;

	component nios_system_rsp_xbar_mux is
		port (
			clk                 : in  std_logic                      := 'X';             -- clk
			reset               : in  std_logic                      := 'X';             -- reset
			src_ready           : in  std_logic                      := 'X';             -- ready
			src_valid           : out std_logic;                                         -- valid
			src_data            : out std_logic_vector(101 downto 0);                    -- data
			src_channel         : out std_logic_vector(7 downto 0);                      -- channel
			src_startofpacket   : out std_logic;                                         -- startofpacket
			src_endofpacket     : out std_logic;                                         -- endofpacket
			sink0_ready         : out std_logic;                                         -- ready
			sink0_valid         : in  std_logic                      := 'X';             -- valid
			sink0_channel       : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- channel
			sink0_data          : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink0_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink0_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink1_ready         : out std_logic;                                         -- ready
			sink1_valid         : in  std_logic                      := 'X';             -- valid
			sink1_channel       : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- channel
			sink1_data          : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink1_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink1_endofpacket   : in  std_logic                      := 'X'              -- endofpacket
		);
	end component nios_system_rsp_xbar_mux;

	component nios_system_rsp_xbar_mux_001 is
		port (
			clk                 : in  std_logic                      := 'X';             -- clk
			reset               : in  std_logic                      := 'X';             -- reset
			src_ready           : in  std_logic                      := 'X';             -- ready
			src_valid           : out std_logic;                                         -- valid
			src_data            : out std_logic_vector(101 downto 0);                    -- data
			src_channel         : out std_logic_vector(7 downto 0);                      -- channel
			src_startofpacket   : out std_logic;                                         -- startofpacket
			src_endofpacket     : out std_logic;                                         -- endofpacket
			sink0_ready         : out std_logic;                                         -- ready
			sink0_valid         : in  std_logic                      := 'X';             -- valid
			sink0_channel       : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- channel
			sink0_data          : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink0_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink0_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink1_ready         : out std_logic;                                         -- ready
			sink1_valid         : in  std_logic                      := 'X';             -- valid
			sink1_channel       : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- channel
			sink1_data          : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink1_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink1_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink2_ready         : out std_logic;                                         -- ready
			sink2_valid         : in  std_logic                      := 'X';             -- valid
			sink2_channel       : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- channel
			sink2_data          : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink2_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink2_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink3_ready         : out std_logic;                                         -- ready
			sink3_valid         : in  std_logic                      := 'X';             -- valid
			sink3_channel       : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- channel
			sink3_data          : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink3_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink3_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink4_ready         : out std_logic;                                         -- ready
			sink4_valid         : in  std_logic                      := 'X';             -- valid
			sink4_channel       : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- channel
			sink4_data          : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink4_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink4_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink5_ready         : out std_logic;                                         -- ready
			sink5_valid         : in  std_logic                      := 'X';             -- valid
			sink5_channel       : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- channel
			sink5_data          : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink5_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink5_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink6_ready         : out std_logic;                                         -- ready
			sink6_valid         : in  std_logic                      := 'X';             -- valid
			sink6_channel       : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- channel
			sink6_data          : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink6_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink6_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink7_ready         : out std_logic;                                         -- ready
			sink7_valid         : in  std_logic                      := 'X';             -- valid
			sink7_channel       : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- channel
			sink7_data          : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink7_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink7_endofpacket   : in  std_logic                      := 'X'              -- endofpacket
		);
	end component nios_system_rsp_xbar_mux_001;

	component nios_system_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component nios_system_irq_mapper;

	component nios_system_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo is
		generic (
			SYMBOLS_PER_BEAT    : integer := 1;
			BITS_PER_SYMBOL     : integer := 8;
			FIFO_DEPTH          : integer := 16;
			CHANNEL_WIDTH       : integer := 0;
			ERROR_WIDTH         : integer := 0;
			USE_PACKETS         : integer := 0;
			USE_FILL_LEVEL      : integer := 0;
			EMPTY_LATENCY       : integer := 3;
			USE_MEMORY_BLOCKS   : integer := 1;
			USE_STORE_FORWARD   : integer := 0;
			USE_ALMOST_FULL_IF  : integer := 0;
			USE_ALMOST_EMPTY_IF : integer := 0
		);
		port (
			clk               : in  std_logic                      := 'X';             -- clk
			reset             : in  std_logic                      := 'X';             -- reset
			in_data           : in  std_logic_vector(102 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                      := 'X';             -- valid
			in_ready          : out std_logic;                                         -- ready
			in_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			out_data          : out std_logic_vector(102 downto 0);                    -- data
			out_valid         : out std_logic;                                         -- valid
			out_ready         : in  std_logic                      := 'X';             -- ready
			out_startofpacket : out std_logic;                                         -- startofpacket
			out_endofpacket   : out std_logic;                                         -- endofpacket
			csr_address       : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- address
			csr_read          : in  std_logic                      := 'X';             -- read
			csr_write         : in  std_logic                      := 'X';             -- write
			csr_readdata      : out std_logic_vector(31 downto 0);                     -- readdata
			csr_writedata     : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			almost_full_data  : out std_logic;                                         -- data
			almost_empty_data : out std_logic;                                         -- data
			in_empty          : in  std_logic                      := 'X';             -- empty
			out_empty         : out std_logic;                                         -- empty
			in_error          : in  std_logic                      := 'X';             -- error
			out_error         : out std_logic;                                         -- error
			in_channel        : in  std_logic                      := 'X';             -- channel
			out_channel       : out std_logic                                          -- channel
		);
	end component nios_system_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo;

	component nios_system_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo is
		generic (
			SYMBOLS_PER_BEAT    : integer := 1;
			BITS_PER_SYMBOL     : integer := 8;
			FIFO_DEPTH          : integer := 16;
			CHANNEL_WIDTH       : integer := 0;
			ERROR_WIDTH         : integer := 0;
			USE_PACKETS         : integer := 0;
			USE_FILL_LEVEL      : integer := 0;
			EMPTY_LATENCY       : integer := 3;
			USE_MEMORY_BLOCKS   : integer := 1;
			USE_STORE_FORWARD   : integer := 0;
			USE_ALMOST_FULL_IF  : integer := 0;
			USE_ALMOST_EMPTY_IF : integer := 0
		);
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			in_data           : in  std_logic_vector(84 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                     := 'X';             -- valid
			in_ready          : out std_logic;                                        -- ready
			in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			out_data          : out std_logic_vector(84 downto 0);                    -- data
			out_valid         : out std_logic;                                        -- valid
			out_ready         : in  std_logic                     := 'X';             -- ready
			out_startofpacket : out std_logic;                                        -- startofpacket
			out_endofpacket   : out std_logic;                                        -- endofpacket
			csr_address       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			csr_read          : in  std_logic                     := 'X';             -- read
			csr_write         : in  std_logic                     := 'X';             -- write
			csr_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			csr_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			almost_full_data  : out std_logic;                                        -- data
			almost_empty_data : out std_logic;                                        -- data
			in_empty          : in  std_logic                     := 'X';             -- empty
			out_empty         : out std_logic;                                        -- empty
			in_error          : in  std_logic                     := 'X';             -- error
			out_error         : out std_logic;                                        -- error
			in_channel        : in  std_logic                     := 'X';             -- channel
			out_channel       : out std_logic                                         -- channel
		);
	end component nios_system_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo;

	component nios_system_sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo is
		generic (
			SYMBOLS_PER_BEAT    : integer := 1;
			BITS_PER_SYMBOL     : integer := 8;
			FIFO_DEPTH          : integer := 16;
			CHANNEL_WIDTH       : integer := 0;
			ERROR_WIDTH         : integer := 0;
			USE_PACKETS         : integer := 0;
			USE_FILL_LEVEL      : integer := 0;
			EMPTY_LATENCY       : integer := 3;
			USE_MEMORY_BLOCKS   : integer := 1;
			USE_STORE_FORWARD   : integer := 0;
			USE_ALMOST_FULL_IF  : integer := 0;
			USE_ALMOST_EMPTY_IF : integer := 0
		);
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			in_data           : in  std_logic_vector(17 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                     := 'X';             -- valid
			in_ready          : out std_logic;                                        -- ready
			out_data          : out std_logic_vector(17 downto 0);                    -- data
			out_valid         : out std_logic;                                        -- valid
			out_ready         : in  std_logic                     := 'X';             -- ready
			csr_address       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			csr_read          : in  std_logic                     := 'X';             -- read
			csr_write         : in  std_logic                     := 'X';             -- write
			csr_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			csr_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			almost_full_data  : out std_logic;                                        -- data
			almost_empty_data : out std_logic;                                        -- data
			in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			out_startofpacket : out std_logic;                                        -- startofpacket
			out_endofpacket   : out std_logic;                                        -- endofpacket
			in_empty          : in  std_logic                     := 'X';             -- empty
			out_empty         : out std_logic;                                        -- empty
			in_error          : in  std_logic                     := 'X';             -- error
			out_error         : out std_logic;                                        -- error
			in_channel        : in  std_logic                     := 'X';             -- channel
			out_channel       : out std_logic                                         -- channel
		);
	end component nios_system_sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo;

	component nios_system_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent is
		generic (
			PKT_DATA_H                : integer := 31;
			PKT_DATA_L                : integer := 0;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_SYMBOL_W              : integer := 8;
			PKT_BYTEEN_H              : integer := 71;
			PKT_BYTEEN_L              : integer := 68;
			PKT_ADDR_H                : integer := 63;
			PKT_ADDR_L                : integer := 32;
			PKT_TRANS_COMPRESSED_READ : integer := 67;
			PKT_TRANS_POSTED          : integer := 66;
			PKT_TRANS_WRITE           : integer := 65;
			PKT_TRANS_READ            : integer := 64;
			PKT_TRANS_LOCK            : integer := 87;
			PKT_SRC_ID_H              : integer := 74;
			PKT_SRC_ID_L              : integer := 72;
			PKT_DEST_ID_H             : integer := 77;
			PKT_DEST_ID_L             : integer := 75;
			PKT_BURSTWRAP_H           : integer := 85;
			PKT_BURSTWRAP_L           : integer := 82;
			PKT_BYTE_CNT_H            : integer := 81;
			PKT_BYTE_CNT_L            : integer := 78;
			PKT_PROTECTION_H          : integer := 86;
			PKT_PROTECTION_L          : integer := 86;
			PKT_RESPONSE_STATUS_H     : integer := 89;
			PKT_RESPONSE_STATUS_L     : integer := 88;
			PKT_BURST_SIZE_H          : integer := 92;
			PKT_BURST_SIZE_L          : integer := 90;
			ST_CHANNEL_W              : integer := 8;
			ST_DATA_W                 : integer := 93;
			AVS_BURSTCOUNT_W          : integer := 4;
			SUPPRESS_0_BYTEEN_CMD     : integer := 1;
			PREVENT_FIFO_OVERFLOW     : integer := 0;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                      := 'X';             -- clk
			reset                   : in  std_logic                      := 'X';             -- reset
			m0_address              : out std_logic_vector(28 downto 0);                     -- address
			m0_burstcount           : out std_logic_vector(2 downto 0);                      -- burstcount
			m0_byteenable           : out std_logic_vector(3 downto 0);                      -- byteenable
			m0_debugaccess          : out std_logic;                                         -- debugaccess
			m0_lock                 : out std_logic;                                         -- lock
			m0_readdata             : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                      := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                         -- read
			m0_waitrequest          : in  std_logic                      := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(31 downto 0);                     -- writedata
			m0_write                : out std_logic;                                         -- write
			rp_endofpacket          : out std_logic;                                         -- endofpacket
			rp_ready                : in  std_logic                      := 'X';             -- ready
			rp_valid                : out std_logic;                                         -- valid
			rp_data                 : out std_logic_vector(101 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                         -- startofpacket
			cp_ready                : out std_logic;                                         -- ready
			cp_valid                : in  std_logic                      := 'X';             -- valid
			cp_data                 : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                      := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                      := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                         -- ready
			rf_sink_valid           : in  std_logic                      := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                      := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                      := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(102 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                      := 'X';             -- ready
			rf_source_valid         : out std_logic;                                         -- valid
			rf_source_startofpacket : out std_logic;                                         -- startofpacket
			rf_source_endofpacket   : out std_logic;                                         -- endofpacket
			rf_source_data          : out std_logic_vector(102 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                         -- ready
			rdata_fifo_sink_valid   : in  std_logic                      := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(33 downto 0)  := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                      := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                         -- valid
			rdata_fifo_src_data     : out std_logic_vector(33 downto 0);                     -- data
			m0_response             : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- response
			m0_writeresponserequest : out std_logic;                                         -- writeresponserequest
			m0_writeresponsevalid   : in  std_logic                      := 'X'              -- writeresponsevalid
		);
	end component nios_system_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent;

	component nios_system_sdram_s1_translator_avalon_universal_slave_0_agent is
		generic (
			PKT_DATA_H                : integer := 31;
			PKT_DATA_L                : integer := 0;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_SYMBOL_W              : integer := 8;
			PKT_BYTEEN_H              : integer := 71;
			PKT_BYTEEN_L              : integer := 68;
			PKT_ADDR_H                : integer := 63;
			PKT_ADDR_L                : integer := 32;
			PKT_TRANS_COMPRESSED_READ : integer := 67;
			PKT_TRANS_POSTED          : integer := 66;
			PKT_TRANS_WRITE           : integer := 65;
			PKT_TRANS_READ            : integer := 64;
			PKT_TRANS_LOCK            : integer := 87;
			PKT_SRC_ID_H              : integer := 74;
			PKT_SRC_ID_L              : integer := 72;
			PKT_DEST_ID_H             : integer := 77;
			PKT_DEST_ID_L             : integer := 75;
			PKT_BURSTWRAP_H           : integer := 85;
			PKT_BURSTWRAP_L           : integer := 82;
			PKT_BYTE_CNT_H            : integer := 81;
			PKT_BYTE_CNT_L            : integer := 78;
			PKT_PROTECTION_H          : integer := 86;
			PKT_PROTECTION_L          : integer := 86;
			PKT_RESPONSE_STATUS_H     : integer := 89;
			PKT_RESPONSE_STATUS_L     : integer := 88;
			PKT_BURST_SIZE_H          : integer := 92;
			PKT_BURST_SIZE_L          : integer := 90;
			ST_CHANNEL_W              : integer := 8;
			ST_DATA_W                 : integer := 93;
			AVS_BURSTCOUNT_W          : integer := 4;
			SUPPRESS_0_BYTEEN_CMD     : integer := 1;
			PREVENT_FIFO_OVERFLOW     : integer := 0;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			m0_address              : out std_logic_vector(28 downto 0);                    -- address
			m0_burstcount           : out std_logic_vector(1 downto 0);                     -- burstcount
			m0_byteenable           : out std_logic_vector(1 downto 0);                     -- byteenable
			m0_debugaccess          : out std_logic;                                        -- debugaccess
			m0_lock                 : out std_logic;                                        -- lock
			m0_readdata             : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                        -- read
			m0_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(15 downto 0);                    -- writedata
			m0_write                : out std_logic;                                        -- write
			rp_endofpacket          : out std_logic;                                        -- endofpacket
			rp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : out std_logic;                                        -- valid
			rp_data                 : out std_logic_vector(83 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_ready                : out std_logic;                                        -- ready
			cp_valid                : in  std_logic                     := 'X';             -- valid
			cp_data                 : in  std_logic_vector(83 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                        -- ready
			rf_sink_valid           : in  std_logic                     := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(84 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                     := 'X';             -- ready
			rf_source_valid         : out std_logic;                                        -- valid
			rf_source_startofpacket : out std_logic;                                        -- startofpacket
			rf_source_endofpacket   : out std_logic;                                        -- endofpacket
			rf_source_data          : out std_logic_vector(84 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                        -- ready
			rdata_fifo_sink_valid   : in  std_logic                     := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(17 downto 0) := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                     := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                        -- valid
			rdata_fifo_src_data     : out std_logic_vector(17 downto 0);                    -- data
			m0_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			m0_writeresponserequest : out std_logic;                                        -- writeresponserequest
			m0_writeresponsevalid   : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component nios_system_sdram_s1_translator_avalon_universal_slave_0_agent;

	component nios_system_width_adapter is
		generic (
			IN_PKT_ADDR_H                 : integer := 60;
			IN_PKT_ADDR_L                 : integer := 36;
			IN_PKT_DATA_H                 : integer := 31;
			IN_PKT_DATA_L                 : integer := 0;
			IN_PKT_BYTEEN_H               : integer := 35;
			IN_PKT_BYTEEN_L               : integer := 32;
			IN_PKT_BYTE_CNT_H             : integer := 63;
			IN_PKT_BYTE_CNT_L             : integer := 61;
			IN_PKT_TRANS_COMPRESSED_READ  : integer := 65;
			IN_PKT_BURSTWRAP_H            : integer := 67;
			IN_PKT_BURSTWRAP_L            : integer := 66;
			IN_PKT_BURST_SIZE_H           : integer := 70;
			IN_PKT_BURST_SIZE_L           : integer := 68;
			IN_PKT_RESPONSE_STATUS_H      : integer := 72;
			IN_PKT_RESPONSE_STATUS_L      : integer := 71;
			IN_PKT_TRANS_EXCLUSIVE        : integer := 73;
			IN_PKT_BURST_TYPE_H           : integer := 75;
			IN_PKT_BURST_TYPE_L           : integer := 74;
			IN_ST_DATA_W                  : integer := 76;
			OUT_PKT_ADDR_H                : integer := 60;
			OUT_PKT_ADDR_L                : integer := 36;
			OUT_PKT_DATA_H                : integer := 31;
			OUT_PKT_DATA_L                : integer := 0;
			OUT_PKT_BYTEEN_H              : integer := 35;
			OUT_PKT_BYTEEN_L              : integer := 32;
			OUT_PKT_BYTE_CNT_H            : integer := 63;
			OUT_PKT_BYTE_CNT_L            : integer := 61;
			OUT_PKT_TRANS_COMPRESSED_READ : integer := 65;
			OUT_PKT_BURST_SIZE_H          : integer := 68;
			OUT_PKT_BURST_SIZE_L          : integer := 66;
			OUT_PKT_RESPONSE_STATUS_H     : integer := 70;
			OUT_PKT_RESPONSE_STATUS_L     : integer := 69;
			OUT_PKT_TRANS_EXCLUSIVE       : integer := 71;
			OUT_PKT_BURST_TYPE_H          : integer := 73;
			OUT_PKT_BURST_TYPE_L          : integer := 72;
			OUT_ST_DATA_W                 : integer := 74;
			ST_CHANNEL_W                  : integer := 32;
			OPTIMIZE_FOR_RSP              : integer := 0;
			RESPONSE_PATH                 : integer := 0
		);
		port (
			clk                  : in  std_logic                      := 'X';             -- clk
			reset                : in  std_logic                      := 'X';             -- reset
			in_valid             : in  std_logic                      := 'X';             -- valid
			in_channel           : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- channel
			in_startofpacket     : in  std_logic                      := 'X';             -- startofpacket
			in_endofpacket       : in  std_logic                      := 'X';             -- endofpacket
			in_ready             : out std_logic;                                         -- ready
			in_data              : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			out_endofpacket      : out std_logic;                                         -- endofpacket
			out_data             : out std_logic_vector(83 downto 0);                     -- data
			out_channel          : out std_logic_vector(7 downto 0);                      -- channel
			out_valid            : out std_logic;                                         -- valid
			out_ready            : in  std_logic                      := 'X';             -- ready
			out_startofpacket    : out std_logic;                                         -- startofpacket
			in_command_size_data : in  std_logic_vector(2 downto 0)   := (others => 'X')  -- data
		);
	end component nios_system_width_adapter;

	component nios_system_width_adapter_001 is
		generic (
			IN_PKT_ADDR_H                 : integer := 60;
			IN_PKT_ADDR_L                 : integer := 36;
			IN_PKT_DATA_H                 : integer := 31;
			IN_PKT_DATA_L                 : integer := 0;
			IN_PKT_BYTEEN_H               : integer := 35;
			IN_PKT_BYTEEN_L               : integer := 32;
			IN_PKT_BYTE_CNT_H             : integer := 63;
			IN_PKT_BYTE_CNT_L             : integer := 61;
			IN_PKT_TRANS_COMPRESSED_READ  : integer := 65;
			IN_PKT_BURSTWRAP_H            : integer := 67;
			IN_PKT_BURSTWRAP_L            : integer := 66;
			IN_PKT_BURST_SIZE_H           : integer := 70;
			IN_PKT_BURST_SIZE_L           : integer := 68;
			IN_PKT_RESPONSE_STATUS_H      : integer := 72;
			IN_PKT_RESPONSE_STATUS_L      : integer := 71;
			IN_PKT_TRANS_EXCLUSIVE        : integer := 73;
			IN_PKT_BURST_TYPE_H           : integer := 75;
			IN_PKT_BURST_TYPE_L           : integer := 74;
			IN_ST_DATA_W                  : integer := 76;
			OUT_PKT_ADDR_H                : integer := 60;
			OUT_PKT_ADDR_L                : integer := 36;
			OUT_PKT_DATA_H                : integer := 31;
			OUT_PKT_DATA_L                : integer := 0;
			OUT_PKT_BYTEEN_H              : integer := 35;
			OUT_PKT_BYTEEN_L              : integer := 32;
			OUT_PKT_BYTE_CNT_H            : integer := 63;
			OUT_PKT_BYTE_CNT_L            : integer := 61;
			OUT_PKT_TRANS_COMPRESSED_READ : integer := 65;
			OUT_PKT_BURST_SIZE_H          : integer := 68;
			OUT_PKT_BURST_SIZE_L          : integer := 66;
			OUT_PKT_RESPONSE_STATUS_H     : integer := 70;
			OUT_PKT_RESPONSE_STATUS_L     : integer := 69;
			OUT_PKT_TRANS_EXCLUSIVE       : integer := 71;
			OUT_PKT_BURST_TYPE_H          : integer := 73;
			OUT_PKT_BURST_TYPE_L          : integer := 72;
			OUT_ST_DATA_W                 : integer := 74;
			ST_CHANNEL_W                  : integer := 32;
			OPTIMIZE_FOR_RSP              : integer := 0;
			RESPONSE_PATH                 : integer := 0
		);
		port (
			clk                  : in  std_logic                      := 'X';             -- clk
			reset                : in  std_logic                      := 'X';             -- reset
			in_valid             : in  std_logic                      := 'X';             -- valid
			in_channel           : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- channel
			in_startofpacket     : in  std_logic                      := 'X';             -- startofpacket
			in_endofpacket       : in  std_logic                      := 'X';             -- endofpacket
			in_ready             : out std_logic;                                         -- ready
			in_data              : in  std_logic_vector(83 downto 0)  := (others => 'X'); -- data
			out_endofpacket      : out std_logic;                                         -- endofpacket
			out_data             : out std_logic_vector(101 downto 0);                    -- data
			out_channel          : out std_logic_vector(7 downto 0);                      -- channel
			out_valid            : out std_logic;                                         -- valid
			out_ready            : in  std_logic                      := 'X';             -- ready
			out_startofpacket    : out std_logic;                                         -- startofpacket
			in_command_size_data : in  std_logic_vector(2 downto 0)   := (others => 'X')  -- data
		);
	end component nios_system_width_adapter_001;

	component nios_system_cpu_instruction_master_translator is
		generic (
			AV_ADDRESS_W                : integer := 32;
			AV_DATA_W                   : integer := 32;
			AV_BURSTCOUNT_W             : integer := 4;
			AV_BYTEENABLE_W             : integer := 4;
			UAV_ADDRESS_W               : integer := 38;
			UAV_BURSTCOUNT_W            : integer := 10;
			USE_READ                    : integer := 1;
			USE_WRITE                   : integer := 1;
			USE_BEGINBURSTTRANSFER      : integer := 0;
			USE_BEGINTRANSFER           : integer := 0;
			USE_CHIPSELECT              : integer := 0;
			USE_BURSTCOUNT              : integer := 1;
			USE_READDATAVALID           : integer := 1;
			USE_WAITREQUEST             : integer := 1;
			USE_READRESPONSE            : integer := 0;
			USE_WRITERESPONSE           : integer := 0;
			AV_SYMBOLS_PER_WORD         : integer := 4;
			AV_ADDRESS_SYMBOLS          : integer := 0;
			AV_BURSTCOUNT_SYMBOLS       : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR  : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR : integer := 0;
			AV_LINEWRAPBURSTS           : integer := 0;
			AV_REGISTERINCOMINGSIGNALS  : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : out std_logic_vector(28 downto 0);                    -- address
			uav_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			uav_read                 : out std_logic;                                        -- read
			uav_write                : out std_logic;                                        -- write
			uav_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			uav_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uav_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			uav_lock                 : out std_logic;                                        -- lock
			uav_debugaccess          : out std_logic;                                        -- debugaccess
			av_address               : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			av_waitrequest           : out std_logic;                                        -- waitrequest
			av_read                  : in  std_logic                     := 'X';             -- read
			av_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			av_readdatavalid         : out std_logic;                                        -- readdatavalid
			av_burstcount            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			av_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_beginbursttransfer    : in  std_logic                     := 'X';             -- beginbursttransfer
			av_begintransfer         : in  std_logic                     := 'X';             -- begintransfer
			av_chipselect            : in  std_logic                     := 'X';             -- chipselect
			av_write                 : in  std_logic                     := 'X';             -- write
			av_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_lock                  : in  std_logic                     := 'X';             -- lock
			av_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			uav_clken                : out std_logic;                                        -- clken
			av_clken                 : in  std_logic                     := 'X';             -- clken
			uav_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			av_response              : out std_logic_vector(1 downto 0);                     -- response
			uav_writeresponserequest : out std_logic;                                        -- writeresponserequest
			uav_writeresponsevalid   : in  std_logic                     := 'X';             -- writeresponsevalid
			av_writeresponserequest  : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid    : out std_logic                                         -- writeresponsevalid
		);
	end component nios_system_cpu_instruction_master_translator;

	component nios_system_cpu_data_master_translator is
		generic (
			AV_ADDRESS_W                : integer := 32;
			AV_DATA_W                   : integer := 32;
			AV_BURSTCOUNT_W             : integer := 4;
			AV_BYTEENABLE_W             : integer := 4;
			UAV_ADDRESS_W               : integer := 38;
			UAV_BURSTCOUNT_W            : integer := 10;
			USE_READ                    : integer := 1;
			USE_WRITE                   : integer := 1;
			USE_BEGINBURSTTRANSFER      : integer := 0;
			USE_BEGINTRANSFER           : integer := 0;
			USE_CHIPSELECT              : integer := 0;
			USE_BURSTCOUNT              : integer := 1;
			USE_READDATAVALID           : integer := 1;
			USE_WAITREQUEST             : integer := 1;
			USE_READRESPONSE            : integer := 0;
			USE_WRITERESPONSE           : integer := 0;
			AV_SYMBOLS_PER_WORD         : integer := 4;
			AV_ADDRESS_SYMBOLS          : integer := 0;
			AV_BURSTCOUNT_SYMBOLS       : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR  : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR : integer := 0;
			AV_LINEWRAPBURSTS           : integer := 0;
			AV_REGISTERINCOMINGSIGNALS  : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : out std_logic_vector(28 downto 0);                    -- address
			uav_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			uav_read                 : out std_logic;                                        -- read
			uav_write                : out std_logic;                                        -- write
			uav_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			uav_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uav_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			uav_lock                 : out std_logic;                                        -- lock
			uav_debugaccess          : out std_logic;                                        -- debugaccess
			av_address               : in  std_logic_vector(28 downto 0) := (others => 'X'); -- address
			av_waitrequest           : out std_logic;                                        -- waitrequest
			av_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_read                  : in  std_logic                     := 'X';             -- read
			av_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			av_write                 : in  std_logic                     := 'X';             -- write
			av_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			av_burstcount            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			av_beginbursttransfer    : in  std_logic                     := 'X';             -- beginbursttransfer
			av_begintransfer         : in  std_logic                     := 'X';             -- begintransfer
			av_chipselect            : in  std_logic                     := 'X';             -- chipselect
			av_readdatavalid         : out std_logic;                                        -- readdatavalid
			av_lock                  : in  std_logic                     := 'X';             -- lock
			uav_clken                : out std_logic;                                        -- clken
			av_clken                 : in  std_logic                     := 'X';             -- clken
			uav_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			av_response              : out std_logic_vector(1 downto 0);                     -- response
			uav_writeresponserequest : out std_logic;                                        -- writeresponserequest
			uav_writeresponsevalid   : in  std_logic                     := 'X';             -- writeresponsevalid
			av_writeresponserequest  : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid    : out std_logic                                         -- writeresponsevalid
		);
	end component nios_system_cpu_data_master_translator;

	component nios_system_cpu_jtag_debug_module_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(28 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(8 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component nios_system_cpu_jtag_debug_module_translator;

	component nios_system_sdram_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(28 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(15 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(23 downto 0);                    -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(15 downto 0);                    -- writedata
			av_byteenable            : out std_logic_vector(1 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_chipselect            : out std_logic;                                        -- chipselect
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_writebyteenable       : out std_logic_vector(1 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component nios_system_sdram_s1_translator;

	component nios_system_interval_timer_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(28 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(2 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_readdata              : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(15 downto 0);                    -- writedata
			av_chipselect            : out std_logic;                                        -- chipselect
			av_read                  : out std_logic;                                        -- read
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component nios_system_interval_timer_s1_translator;

	component nios_system_sysid_control_slave_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(28 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(0 downto 0);                     -- address
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component nios_system_sysid_control_slave_translator;

	component nios_system_jtag_uart_avalon_jtag_slave_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(28 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(0 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_chipselect            : out std_logic;                                        -- chipselect
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component nios_system_jtag_uart_avalon_jtag_slave_translator;

	component nios_system_ctr_moteur_avalon_parallel_port_slave_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(28 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(1 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_chipselect            : out std_logic;                                        -- chipselect
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component nios_system_ctr_moteur_avalon_parallel_port_slave_translator;

	component nios_system_rst_controller is
		generic (
			NUM_RESET_INPUTS        : integer := 6;
			OUTPUT_RESET_SYNC_EDGES : string  := "deassert";
			SYNC_DEPTH              : integer := 2;
			RESET_REQUEST_PRESENT   : integer := 0
		);
		port (
			reset_in0  : in  std_logic := 'X'; -- reset
			reset_in1  : in  std_logic := 'X'; -- reset
			clk        : in  std_logic := 'X'; -- clk
			reset_out  : out std_logic;        -- reset
			reset_req  : out std_logic;        -- reset_req
			reset_in2  : in  std_logic := 'X'; -- reset
			reset_in3  : in  std_logic := 'X'; -- reset
			reset_in4  : in  std_logic := 'X'; -- reset
			reset_in5  : in  std_logic := 'X'; -- reset
			reset_in6  : in  std_logic := 'X'; -- reset
			reset_in7  : in  std_logic := 'X'; -- reset
			reset_in8  : in  std_logic := 'X'; -- reset
			reset_in9  : in  std_logic := 'X'; -- reset
			reset_in10 : in  std_logic := 'X'; -- reset
			reset_in11 : in  std_logic := 'X'; -- reset
			reset_in12 : in  std_logic := 'X'; -- reset
			reset_in13 : in  std_logic := 'X'; -- reset
			reset_in14 : in  std_logic := 'X'; -- reset
			reset_in15 : in  std_logic := 'X'  -- reset
		);
	end component nios_system_rst_controller;

	component nios_system_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS        : integer := 6;
			OUTPUT_RESET_SYNC_EDGES : string  := "deassert";
			SYNC_DEPTH              : integer := 2;
			RESET_REQUEST_PRESENT   : integer := 0
		);
		port (
			reset_in0  : in  std_logic := 'X'; -- reset
			clk        : in  std_logic := 'X'; -- clk
			reset_out  : out std_logic;        -- reset
			reset_req  : out std_logic;        -- reset_req
			reset_in1  : in  std_logic := 'X'; -- reset
			reset_in2  : in  std_logic := 'X'; -- reset
			reset_in3  : in  std_logic := 'X'; -- reset
			reset_in4  : in  std_logic := 'X'; -- reset
			reset_in5  : in  std_logic := 'X'; -- reset
			reset_in6  : in  std_logic := 'X'; -- reset
			reset_in7  : in  std_logic := 'X'; -- reset
			reset_in8  : in  std_logic := 'X'; -- reset
			reset_in9  : in  std_logic := 'X'; -- reset
			reset_in10 : in  std_logic := 'X'; -- reset
			reset_in11 : in  std_logic := 'X'; -- reset
			reset_in12 : in  std_logic := 'X'; -- reset
			reset_in13 : in  std_logic := 'X'; -- reset
			reset_in14 : in  std_logic := 'X'; -- reset
			reset_in15 : in  std_logic := 'X'  -- reset
		);
	end component nios_system_rst_controller_001;

	signal external_clocks_sys_clk_clk                                                                                : std_logic;                      -- External_Clocks:sys_clk -> [CPU:clk, CPU_data_master_translator:clk, CPU_data_master_translator_avalon_universal_master_0_agent:clk, CPU_instruction_master_translator:clk, CPU_instruction_master_translator_avalon_universal_master_0_agent:clk, CPU_jtag_debug_module_translator:clk, CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:clk, CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, CTR_MOTEUR:clk, CTR_MOTEUR_avalon_parallel_port_slave_translator:clk, CTR_MOTEUR_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:clk, CTR_MOTEUR_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Interval_timer:clk, Interval_timer_s1_translator:clk, Interval_timer_s1_translator_avalon_universal_slave_0_agent:clk, Interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, JTAG_UART:clk, JTAG_UART_avalon_jtag_slave_translator:clk, JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:clk, JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, SDRAM:clk, SDRAM_s1_translator:clk, SDRAM_s1_translator_avalon_universal_slave_0_agent:clk, SDRAM_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, SDRAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, addr_router:clk, addr_router_001:clk, burst_adapter:clk, capt3_0:clk, capt3_0_avalon_parallel_port_slave_translator:clk, capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:clk, capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, capt6_4:clk, capt6_4_avalon_parallel_port_slave_translator:clk, capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:clk, capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, cmd_xbar_demux:clk, cmd_xbar_demux_001:clk, cmd_xbar_mux:clk, cmd_xbar_mux_001:clk, id_router:clk, id_router_001:clk, id_router_002:clk, id_router_003:clk, id_router_004:clk, id_router_005:clk, id_router_006:clk, id_router_007:clk, irq_mapper:clk, limiter:clk, rsp_xbar_demux:clk, rsp_xbar_demux_001:clk, rsp_xbar_demux_002:clk, rsp_xbar_demux_003:clk, rsp_xbar_demux_004:clk, rsp_xbar_demux_005:clk, rsp_xbar_demux_006:clk, rsp_xbar_demux_007:clk, rsp_xbar_mux:clk, rsp_xbar_mux_001:clk, rst_controller:clk, sysid:clock, sysid_control_slave_translator:clk, sysid_control_slave_translator_avalon_universal_slave_0_agent:clk, sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, width_adapter:clk, width_adapter_001:clk]
	signal cpu_jtag_debug_module_reset_reset                                                                          : std_logic;                      -- CPU:jtag_debug_module_resetrequest -> [CTR_MOTEUR:reset, CTR_MOTEUR_avalon_parallel_port_slave_translator:reset, CTR_MOTEUR_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:reset, CTR_MOTEUR_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, capt3_0:reset, capt3_0_avalon_parallel_port_slave_translator:reset, capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:reset, capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, capt6_4:reset, capt6_4_avalon_parallel_port_slave_translator:reset, capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:reset, capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router_005:reset, id_router_006:reset, id_router_007:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rst_controller:reset_in1]
	signal cpu_instruction_master_waitrequest                                                                         : std_logic;                      -- CPU_instruction_master_translator:av_waitrequest -> CPU:i_waitrequest
	signal cpu_instruction_master_address                                                                             : std_logic_vector(27 downto 0);  -- CPU:i_address -> CPU_instruction_master_translator:av_address
	signal cpu_instruction_master_read                                                                                : std_logic;                      -- CPU:i_read -> CPU_instruction_master_translator:av_read
	signal cpu_instruction_master_readdata                                                                            : std_logic_vector(31 downto 0);  -- CPU_instruction_master_translator:av_readdata -> CPU:i_readdata
	signal cpu_instruction_master_readdatavalid                                                                       : std_logic;                      -- CPU_instruction_master_translator:av_readdatavalid -> CPU:i_readdatavalid
	signal cpu_data_master_waitrequest                                                                                : std_logic;                      -- CPU_data_master_translator:av_waitrequest -> CPU:d_waitrequest
	signal cpu_data_master_writedata                                                                                  : std_logic_vector(31 downto 0);  -- CPU:d_writedata -> CPU_data_master_translator:av_writedata
	signal cpu_data_master_address                                                                                    : std_logic_vector(28 downto 0);  -- CPU:d_address -> CPU_data_master_translator:av_address
	signal cpu_data_master_write                                                                                      : std_logic;                      -- CPU:d_write -> CPU_data_master_translator:av_write
	signal cpu_data_master_read                                                                                       : std_logic;                      -- CPU:d_read -> CPU_data_master_translator:av_read
	signal cpu_data_master_readdata                                                                                   : std_logic_vector(31 downto 0);  -- CPU_data_master_translator:av_readdata -> CPU:d_readdata
	signal cpu_data_master_debugaccess                                                                                : std_logic;                      -- CPU:jtag_debug_module_debugaccess_to_roms -> CPU_data_master_translator:av_debugaccess
	signal cpu_data_master_byteenable                                                                                 : std_logic_vector(3 downto 0);   -- CPU:d_byteenable -> CPU_data_master_translator:av_byteenable
	signal cpu_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest                                           : std_logic;                      -- CPU:jtag_debug_module_waitrequest -> CPU_jtag_debug_module_translator:av_waitrequest
	signal cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata                                             : std_logic_vector(31 downto 0);  -- CPU_jtag_debug_module_translator:av_writedata -> CPU:jtag_debug_module_writedata
	signal cpu_jtag_debug_module_translator_avalon_anti_slave_0_address                                               : std_logic_vector(8 downto 0);   -- CPU_jtag_debug_module_translator:av_address -> CPU:jtag_debug_module_address
	signal cpu_jtag_debug_module_translator_avalon_anti_slave_0_write                                                 : std_logic;                      -- CPU_jtag_debug_module_translator:av_write -> CPU:jtag_debug_module_write
	signal cpu_jtag_debug_module_translator_avalon_anti_slave_0_read                                                  : std_logic;                      -- CPU_jtag_debug_module_translator:av_read -> CPU:jtag_debug_module_read
	signal cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata                                              : std_logic_vector(31 downto 0);  -- CPU:jtag_debug_module_readdata -> CPU_jtag_debug_module_translator:av_readdata
	signal cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess                                           : std_logic;                      -- CPU_jtag_debug_module_translator:av_debugaccess -> CPU:jtag_debug_module_debugaccess
	signal cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable                                            : std_logic_vector(3 downto 0);   -- CPU_jtag_debug_module_translator:av_byteenable -> CPU:jtag_debug_module_byteenable
	signal sdram_s1_translator_avalon_anti_slave_0_waitrequest                                                        : std_logic;                      -- SDRAM:za_waitrequest -> SDRAM_s1_translator:av_waitrequest
	signal sdram_s1_translator_avalon_anti_slave_0_writedata                                                          : std_logic_vector(15 downto 0);  -- SDRAM_s1_translator:av_writedata -> SDRAM:az_data
	signal sdram_s1_translator_avalon_anti_slave_0_address                                                            : std_logic_vector(23 downto 0);  -- SDRAM_s1_translator:av_address -> SDRAM:az_addr
	signal sdram_s1_translator_avalon_anti_slave_0_chipselect                                                         : std_logic;                      -- SDRAM_s1_translator:av_chipselect -> SDRAM:az_cs
	signal sdram_s1_translator_avalon_anti_slave_0_write                                                              : std_logic;                      -- SDRAM_s1_translator:av_write -> sdram_s1_translator_avalon_anti_slave_0_write:in
	signal sdram_s1_translator_avalon_anti_slave_0_read                                                               : std_logic;                      -- SDRAM_s1_translator:av_read -> sdram_s1_translator_avalon_anti_slave_0_read:in
	signal sdram_s1_translator_avalon_anti_slave_0_readdata                                                           : std_logic_vector(15 downto 0);  -- SDRAM:za_data -> SDRAM_s1_translator:av_readdata
	signal sdram_s1_translator_avalon_anti_slave_0_readdatavalid                                                      : std_logic;                      -- SDRAM:za_valid -> SDRAM_s1_translator:av_readdatavalid
	signal sdram_s1_translator_avalon_anti_slave_0_byteenable                                                         : std_logic_vector(1 downto 0);   -- SDRAM_s1_translator:av_byteenable -> sdram_s1_translator_avalon_anti_slave_0_byteenable:in
	signal interval_timer_s1_translator_avalon_anti_slave_0_writedata                                                 : std_logic_vector(15 downto 0);  -- Interval_timer_s1_translator:av_writedata -> Interval_timer:writedata
	signal interval_timer_s1_translator_avalon_anti_slave_0_address                                                   : std_logic_vector(2 downto 0);   -- Interval_timer_s1_translator:av_address -> Interval_timer:address
	signal interval_timer_s1_translator_avalon_anti_slave_0_chipselect                                                : std_logic;                      -- Interval_timer_s1_translator:av_chipselect -> Interval_timer:chipselect
	signal interval_timer_s1_translator_avalon_anti_slave_0_write                                                     : std_logic;                      -- Interval_timer_s1_translator:av_write -> interval_timer_s1_translator_avalon_anti_slave_0_write:in
	signal interval_timer_s1_translator_avalon_anti_slave_0_readdata                                                  : std_logic_vector(15 downto 0);  -- Interval_timer:readdata -> Interval_timer_s1_translator:av_readdata
	signal sysid_control_slave_translator_avalon_anti_slave_0_address                                                 : std_logic_vector(0 downto 0);   -- sysid_control_slave_translator:av_address -> sysid:address
	signal sysid_control_slave_translator_avalon_anti_slave_0_readdata                                                : std_logic_vector(31 downto 0);  -- sysid:readdata -> sysid_control_slave_translator:av_readdata
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest                                     : std_logic;                      -- JTAG_UART:av_waitrequest -> JTAG_UART_avalon_jtag_slave_translator:av_waitrequest
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata                                       : std_logic_vector(31 downto 0);  -- JTAG_UART_avalon_jtag_slave_translator:av_writedata -> JTAG_UART:av_writedata
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address                                         : std_logic_vector(0 downto 0);   -- JTAG_UART_avalon_jtag_slave_translator:av_address -> JTAG_UART:av_address
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect                                      : std_logic;                      -- JTAG_UART_avalon_jtag_slave_translator:av_chipselect -> JTAG_UART:av_chipselect
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write                                           : std_logic;                      -- JTAG_UART_avalon_jtag_slave_translator:av_write -> jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write:in
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read                                            : std_logic;                      -- JTAG_UART_avalon_jtag_slave_translator:av_read -> jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read:in
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata                                        : std_logic_vector(31 downto 0);  -- JTAG_UART:av_readdata -> JTAG_UART_avalon_jtag_slave_translator:av_readdata
	signal ctr_moteur_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata                             : std_logic_vector(31 downto 0);  -- CTR_MOTEUR_avalon_parallel_port_slave_translator:av_writedata -> CTR_MOTEUR:writedata
	signal ctr_moteur_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address                               : std_logic_vector(1 downto 0);   -- CTR_MOTEUR_avalon_parallel_port_slave_translator:av_address -> CTR_MOTEUR:address
	signal ctr_moteur_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect                            : std_logic;                      -- CTR_MOTEUR_avalon_parallel_port_slave_translator:av_chipselect -> CTR_MOTEUR:chipselect
	signal ctr_moteur_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write                                 : std_logic;                      -- CTR_MOTEUR_avalon_parallel_port_slave_translator:av_write -> CTR_MOTEUR:write
	signal ctr_moteur_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read                                  : std_logic;                      -- CTR_MOTEUR_avalon_parallel_port_slave_translator:av_read -> CTR_MOTEUR:read
	signal ctr_moteur_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata                              : std_logic_vector(31 downto 0);  -- CTR_MOTEUR:readdata -> CTR_MOTEUR_avalon_parallel_port_slave_translator:av_readdata
	signal ctr_moteur_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable                            : std_logic_vector(3 downto 0);   -- CTR_MOTEUR_avalon_parallel_port_slave_translator:av_byteenable -> CTR_MOTEUR:byteenable
	signal capt3_0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata                                : std_logic_vector(31 downto 0);  -- capt3_0_avalon_parallel_port_slave_translator:av_writedata -> capt3_0:writedata
	signal capt3_0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address                                  : std_logic_vector(1 downto 0);   -- capt3_0_avalon_parallel_port_slave_translator:av_address -> capt3_0:address
	signal capt3_0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect                               : std_logic;                      -- capt3_0_avalon_parallel_port_slave_translator:av_chipselect -> capt3_0:chipselect
	signal capt3_0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write                                    : std_logic;                      -- capt3_0_avalon_parallel_port_slave_translator:av_write -> capt3_0:write
	signal capt3_0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read                                     : std_logic;                      -- capt3_0_avalon_parallel_port_slave_translator:av_read -> capt3_0:read
	signal capt3_0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata                                 : std_logic_vector(31 downto 0);  -- capt3_0:readdata -> capt3_0_avalon_parallel_port_slave_translator:av_readdata
	signal capt3_0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable                               : std_logic_vector(3 downto 0);   -- capt3_0_avalon_parallel_port_slave_translator:av_byteenable -> capt3_0:byteenable
	signal capt6_4_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata                                : std_logic_vector(31 downto 0);  -- capt6_4_avalon_parallel_port_slave_translator:av_writedata -> capt6_4:writedata
	signal capt6_4_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address                                  : std_logic_vector(1 downto 0);   -- capt6_4_avalon_parallel_port_slave_translator:av_address -> capt6_4:address
	signal capt6_4_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect                               : std_logic;                      -- capt6_4_avalon_parallel_port_slave_translator:av_chipselect -> capt6_4:chipselect
	signal capt6_4_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write                                    : std_logic;                      -- capt6_4_avalon_parallel_port_slave_translator:av_write -> capt6_4:write
	signal capt6_4_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read                                     : std_logic;                      -- capt6_4_avalon_parallel_port_slave_translator:av_read -> capt6_4:read
	signal capt6_4_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata                                 : std_logic_vector(31 downto 0);  -- capt6_4:readdata -> capt6_4_avalon_parallel_port_slave_translator:av_readdata
	signal capt6_4_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable                               : std_logic_vector(3 downto 0);   -- capt6_4_avalon_parallel_port_slave_translator:av_byteenable -> capt6_4:byteenable
	signal cpu_instruction_master_translator_avalon_universal_master_0_waitrequest                                    : std_logic;                      -- CPU_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> CPU_instruction_master_translator:uav_waitrequest
	signal cpu_instruction_master_translator_avalon_universal_master_0_burstcount                                     : std_logic_vector(2 downto 0);   -- CPU_instruction_master_translator:uav_burstcount -> CPU_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	signal cpu_instruction_master_translator_avalon_universal_master_0_writedata                                      : std_logic_vector(31 downto 0);  -- CPU_instruction_master_translator:uav_writedata -> CPU_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	signal cpu_instruction_master_translator_avalon_universal_master_0_address                                        : std_logic_vector(28 downto 0);  -- CPU_instruction_master_translator:uav_address -> CPU_instruction_master_translator_avalon_universal_master_0_agent:av_address
	signal cpu_instruction_master_translator_avalon_universal_master_0_lock                                           : std_logic;                      -- CPU_instruction_master_translator:uav_lock -> CPU_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	signal cpu_instruction_master_translator_avalon_universal_master_0_write                                          : std_logic;                      -- CPU_instruction_master_translator:uav_write -> CPU_instruction_master_translator_avalon_universal_master_0_agent:av_write
	signal cpu_instruction_master_translator_avalon_universal_master_0_read                                           : std_logic;                      -- CPU_instruction_master_translator:uav_read -> CPU_instruction_master_translator_avalon_universal_master_0_agent:av_read
	signal cpu_instruction_master_translator_avalon_universal_master_0_readdata                                       : std_logic_vector(31 downto 0);  -- CPU_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> CPU_instruction_master_translator:uav_readdata
	signal cpu_instruction_master_translator_avalon_universal_master_0_debugaccess                                    : std_logic;                      -- CPU_instruction_master_translator:uav_debugaccess -> CPU_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	signal cpu_instruction_master_translator_avalon_universal_master_0_byteenable                                     : std_logic_vector(3 downto 0);   -- CPU_instruction_master_translator:uav_byteenable -> CPU_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	signal cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid                                  : std_logic;                      -- CPU_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> CPU_instruction_master_translator:uav_readdatavalid
	signal cpu_data_master_translator_avalon_universal_master_0_waitrequest                                           : std_logic;                      -- CPU_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> CPU_data_master_translator:uav_waitrequest
	signal cpu_data_master_translator_avalon_universal_master_0_burstcount                                            : std_logic_vector(2 downto 0);   -- CPU_data_master_translator:uav_burstcount -> CPU_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	signal cpu_data_master_translator_avalon_universal_master_0_writedata                                             : std_logic_vector(31 downto 0);  -- CPU_data_master_translator:uav_writedata -> CPU_data_master_translator_avalon_universal_master_0_agent:av_writedata
	signal cpu_data_master_translator_avalon_universal_master_0_address                                               : std_logic_vector(28 downto 0);  -- CPU_data_master_translator:uav_address -> CPU_data_master_translator_avalon_universal_master_0_agent:av_address
	signal cpu_data_master_translator_avalon_universal_master_0_lock                                                  : std_logic;                      -- CPU_data_master_translator:uav_lock -> CPU_data_master_translator_avalon_universal_master_0_agent:av_lock
	signal cpu_data_master_translator_avalon_universal_master_0_write                                                 : std_logic;                      -- CPU_data_master_translator:uav_write -> CPU_data_master_translator_avalon_universal_master_0_agent:av_write
	signal cpu_data_master_translator_avalon_universal_master_0_read                                                  : std_logic;                      -- CPU_data_master_translator:uav_read -> CPU_data_master_translator_avalon_universal_master_0_agent:av_read
	signal cpu_data_master_translator_avalon_universal_master_0_readdata                                              : std_logic_vector(31 downto 0);  -- CPU_data_master_translator_avalon_universal_master_0_agent:av_readdata -> CPU_data_master_translator:uav_readdata
	signal cpu_data_master_translator_avalon_universal_master_0_debugaccess                                           : std_logic;                      -- CPU_data_master_translator:uav_debugaccess -> CPU_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	signal cpu_data_master_translator_avalon_universal_master_0_byteenable                                            : std_logic_vector(3 downto 0);   -- CPU_data_master_translator:uav_byteenable -> CPU_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	signal cpu_data_master_translator_avalon_universal_master_0_readdatavalid                                         : std_logic;                      -- CPU_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> CPU_data_master_translator:uav_readdatavalid
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest                             : std_logic;                      -- CPU_jtag_debug_module_translator:uav_waitrequest -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount                              : std_logic_vector(2 downto 0);   -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> CPU_jtag_debug_module_translator:uav_burstcount
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata                               : std_logic_vector(31 downto 0);  -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> CPU_jtag_debug_module_translator:uav_writedata
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address                                 : std_logic_vector(28 downto 0);  -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> CPU_jtag_debug_module_translator:uav_address
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write                                   : std_logic;                      -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> CPU_jtag_debug_module_translator:uav_write
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock                                    : std_logic;                      -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> CPU_jtag_debug_module_translator:uav_lock
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read                                    : std_logic;                      -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> CPU_jtag_debug_module_translator:uav_read
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata                                : std_logic_vector(31 downto 0);  -- CPU_jtag_debug_module_translator:uav_readdata -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid                           : std_logic;                      -- CPU_jtag_debug_module_translator:uav_readdatavalid -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess                             : std_logic;                      -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CPU_jtag_debug_module_translator:uav_debugaccess
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable                              : std_logic_vector(3 downto 0);   -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> CPU_jtag_debug_module_translator:uav_byteenable
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                      : std_logic;                      -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid                            : std_logic;                      -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                    : std_logic;                      -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data                             : std_logic_vector(102 downto 0); -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready                            : std_logic;                      -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                   : std_logic;                      -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                         : std_logic;                      -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                 : std_logic;                      -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                          : std_logic_vector(102 downto 0); -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                         : std_logic;                      -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                       : std_logic;                      -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                        : std_logic_vector(33 downto 0);  -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                       : std_logic;                      -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                          : std_logic;                      -- SDRAM_s1_translator:uav_waitrequest -> SDRAM_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                           : std_logic_vector(1 downto 0);   -- SDRAM_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> SDRAM_s1_translator:uav_burstcount
	signal sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                            : std_logic_vector(15 downto 0);  -- SDRAM_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> SDRAM_s1_translator:uav_writedata
	signal sdram_s1_translator_avalon_universal_slave_0_agent_m0_address                                              : std_logic_vector(28 downto 0);  -- SDRAM_s1_translator_avalon_universal_slave_0_agent:m0_address -> SDRAM_s1_translator:uav_address
	signal sdram_s1_translator_avalon_universal_slave_0_agent_m0_write                                                : std_logic;                      -- SDRAM_s1_translator_avalon_universal_slave_0_agent:m0_write -> SDRAM_s1_translator:uav_write
	signal sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock                                                 : std_logic;                      -- SDRAM_s1_translator_avalon_universal_slave_0_agent:m0_lock -> SDRAM_s1_translator:uav_lock
	signal sdram_s1_translator_avalon_universal_slave_0_agent_m0_read                                                 : std_logic;                      -- SDRAM_s1_translator_avalon_universal_slave_0_agent:m0_read -> SDRAM_s1_translator:uav_read
	signal sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                             : std_logic_vector(15 downto 0);  -- SDRAM_s1_translator:uav_readdata -> SDRAM_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                        : std_logic;                      -- SDRAM_s1_translator:uav_readdatavalid -> SDRAM_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                          : std_logic;                      -- SDRAM_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> SDRAM_s1_translator:uav_debugaccess
	signal sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                           : std_logic_vector(1 downto 0);   -- SDRAM_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> SDRAM_s1_translator:uav_byteenable
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                                   : std_logic;                      -- SDRAM_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> SDRAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                         : std_logic;                      -- SDRAM_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> SDRAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                                 : std_logic;                      -- SDRAM_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> SDRAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                          : std_logic_vector(84 downto 0);  -- SDRAM_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> SDRAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                         : std_logic;                      -- SDRAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> SDRAM_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                                : std_logic;                      -- SDRAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> SDRAM_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                      : std_logic;                      -- SDRAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> SDRAM_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                              : std_logic;                      -- SDRAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> SDRAM_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                       : std_logic_vector(84 downto 0);  -- SDRAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> SDRAM_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                      : std_logic;                      -- SDRAM_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> SDRAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                                    : std_logic;                      -- SDRAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> SDRAM_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                                     : std_logic_vector(17 downto 0);  -- SDRAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> SDRAM_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                                    : std_logic;                      -- SDRAM_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> SDRAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid                                    : std_logic;                      -- SDRAM_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> SDRAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data                                     : std_logic_vector(17 downto 0);  -- SDRAM_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> SDRAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready                                    : std_logic;                      -- SDRAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> SDRAM_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	signal interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                 : std_logic;                      -- Interval_timer_s1_translator:uav_waitrequest -> Interval_timer_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                  : std_logic_vector(2 downto 0);   -- Interval_timer_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> Interval_timer_s1_translator:uav_burstcount
	signal interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                   : std_logic_vector(31 downto 0);  -- Interval_timer_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> Interval_timer_s1_translator:uav_writedata
	signal interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_address                                     : std_logic_vector(28 downto 0);  -- Interval_timer_s1_translator_avalon_universal_slave_0_agent:m0_address -> Interval_timer_s1_translator:uav_address
	signal interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_write                                       : std_logic;                      -- Interval_timer_s1_translator_avalon_universal_slave_0_agent:m0_write -> Interval_timer_s1_translator:uav_write
	signal interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock                                        : std_logic;                      -- Interval_timer_s1_translator_avalon_universal_slave_0_agent:m0_lock -> Interval_timer_s1_translator:uav_lock
	signal interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_read                                        : std_logic;                      -- Interval_timer_s1_translator_avalon_universal_slave_0_agent:m0_read -> Interval_timer_s1_translator:uav_read
	signal interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                    : std_logic_vector(31 downto 0);  -- Interval_timer_s1_translator:uav_readdata -> Interval_timer_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                               : std_logic;                      -- Interval_timer_s1_translator:uav_readdatavalid -> Interval_timer_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                 : std_logic;                      -- Interval_timer_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Interval_timer_s1_translator:uav_debugaccess
	signal interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                  : std_logic_vector(3 downto 0);   -- Interval_timer_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> Interval_timer_s1_translator:uav_byteenable
	signal interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                          : std_logic;                      -- Interval_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                : std_logic;                      -- Interval_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> Interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                        : std_logic;                      -- Interval_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                 : std_logic_vector(102 downto 0); -- Interval_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> Interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                : std_logic;                      -- Interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Interval_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                       : std_logic;                      -- Interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Interval_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                             : std_logic;                      -- Interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Interval_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                     : std_logic;                      -- Interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Interval_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                              : std_logic_vector(102 downto 0); -- Interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Interval_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                             : std_logic;                      -- Interval_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal interval_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                           : std_logic;                      -- Interval_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Interval_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal interval_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                            : std_logic_vector(33 downto 0);  -- Interval_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Interval_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal interval_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                           : std_logic;                      -- Interval_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Interval_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest                               : std_logic;                      -- sysid_control_slave_translator:uav_waitrequest -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount                                : std_logic_vector(2 downto 0);   -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> sysid_control_slave_translator:uav_burstcount
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata                                 : std_logic_vector(31 downto 0);  -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> sysid_control_slave_translator:uav_writedata
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address                                   : std_logic_vector(28 downto 0);  -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> sysid_control_slave_translator:uav_address
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write                                     : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> sysid_control_slave_translator:uav_write
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock                                      : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> sysid_control_slave_translator:uav_lock
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read                                      : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> sysid_control_slave_translator:uav_read
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata                                  : std_logic_vector(31 downto 0);  -- sysid_control_slave_translator:uav_readdata -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid                             : std_logic;                      -- sysid_control_slave_translator:uav_readdatavalid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess                               : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sysid_control_slave_translator:uav_debugaccess
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable                                : std_logic_vector(3 downto 0);   -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> sysid_control_slave_translator:uav_byteenable
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                        : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid                              : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                      : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data                               : std_logic_vector(102 downto 0); -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready                              : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                     : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                           : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                   : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                            : std_logic_vector(102 downto 0); -- sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                           : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                         : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                          : std_logic_vector(33 downto 0);  -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                         : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest                       : std_logic;                      -- JTAG_UART_avalon_jtag_slave_translator:uav_waitrequest -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount                        : std_logic_vector(2 downto 0);   -- JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> JTAG_UART_avalon_jtag_slave_translator:uav_burstcount
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata                         : std_logic_vector(31 downto 0);  -- JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> JTAG_UART_avalon_jtag_slave_translator:uav_writedata
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address                           : std_logic_vector(28 downto 0);  -- JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> JTAG_UART_avalon_jtag_slave_translator:uav_address
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write                             : std_logic;                      -- JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> JTAG_UART_avalon_jtag_slave_translator:uav_write
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock                              : std_logic;                      -- JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> JTAG_UART_avalon_jtag_slave_translator:uav_lock
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read                              : std_logic;                      -- JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> JTAG_UART_avalon_jtag_slave_translator:uav_read
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata                          : std_logic_vector(31 downto 0);  -- JTAG_UART_avalon_jtag_slave_translator:uav_readdata -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid                     : std_logic;                      -- JTAG_UART_avalon_jtag_slave_translator:uav_readdatavalid -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess                       : std_logic;                      -- JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> JTAG_UART_avalon_jtag_slave_translator:uav_debugaccess
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable                        : std_logic_vector(3 downto 0);   -- JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> JTAG_UART_avalon_jtag_slave_translator:uav_byteenable
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                : std_logic;                      -- JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid                      : std_logic;                      -- JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket              : std_logic;                      -- JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data                       : std_logic_vector(102 downto 0); -- JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready                      : std_logic;                      -- JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket             : std_logic;                      -- JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                   : std_logic;                      -- JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket           : std_logic;                      -- JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                    : std_logic_vector(102 downto 0); -- JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                   : std_logic;                      -- JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                 : std_logic;                      -- JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                  : std_logic_vector(33 downto 0);  -- JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                 : std_logic;                      -- JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest             : std_logic;                      -- CTR_MOTEUR_avalon_parallel_port_slave_translator:uav_waitrequest -> CTR_MOTEUR_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount              : std_logic_vector(2 downto 0);   -- CTR_MOTEUR_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> CTR_MOTEUR_avalon_parallel_port_slave_translator:uav_burstcount
	signal ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata               : std_logic_vector(31 downto 0);  -- CTR_MOTEUR_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> CTR_MOTEUR_avalon_parallel_port_slave_translator:uav_writedata
	signal ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address                 : std_logic_vector(28 downto 0);  -- CTR_MOTEUR_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_address -> CTR_MOTEUR_avalon_parallel_port_slave_translator:uav_address
	signal ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write                   : std_logic;                      -- CTR_MOTEUR_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_write -> CTR_MOTEUR_avalon_parallel_port_slave_translator:uav_write
	signal ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock                    : std_logic;                      -- CTR_MOTEUR_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_lock -> CTR_MOTEUR_avalon_parallel_port_slave_translator:uav_lock
	signal ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read                    : std_logic;                      -- CTR_MOTEUR_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_read -> CTR_MOTEUR_avalon_parallel_port_slave_translator:uav_read
	signal ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata                : std_logic_vector(31 downto 0);  -- CTR_MOTEUR_avalon_parallel_port_slave_translator:uav_readdata -> CTR_MOTEUR_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid           : std_logic;                      -- CTR_MOTEUR_avalon_parallel_port_slave_translator:uav_readdatavalid -> CTR_MOTEUR_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess             : std_logic;                      -- CTR_MOTEUR_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CTR_MOTEUR_avalon_parallel_port_slave_translator:uav_debugaccess
	signal ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable              : std_logic_vector(3 downto 0);   -- CTR_MOTEUR_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> CTR_MOTEUR_avalon_parallel_port_slave_translator:uav_byteenable
	signal ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket      : std_logic;                      -- CTR_MOTEUR_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CTR_MOTEUR_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid            : std_logic;                      -- CTR_MOTEUR_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> CTR_MOTEUR_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket    : std_logic;                      -- CTR_MOTEUR_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CTR_MOTEUR_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data             : std_logic_vector(102 downto 0); -- CTR_MOTEUR_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> CTR_MOTEUR_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready            : std_logic;                      -- CTR_MOTEUR_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CTR_MOTEUR_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket   : std_logic;                      -- CTR_MOTEUR_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CTR_MOTEUR_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid         : std_logic;                      -- CTR_MOTEUR_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CTR_MOTEUR_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket : std_logic;                      -- CTR_MOTEUR_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CTR_MOTEUR_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data          : std_logic_vector(102 downto 0); -- CTR_MOTEUR_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CTR_MOTEUR_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready         : std_logic;                      -- CTR_MOTEUR_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CTR_MOTEUR_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid       : std_logic;                      -- CTR_MOTEUR_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CTR_MOTEUR_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data        : std_logic_vector(33 downto 0);  -- CTR_MOTEUR_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CTR_MOTEUR_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready       : std_logic;                      -- CTR_MOTEUR_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CTR_MOTEUR_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest                : std_logic;                      -- capt3_0_avalon_parallel_port_slave_translator:uav_waitrequest -> capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount                 : std_logic_vector(2 downto 0);   -- capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> capt3_0_avalon_parallel_port_slave_translator:uav_burstcount
	signal capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata                  : std_logic_vector(31 downto 0);  -- capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> capt3_0_avalon_parallel_port_slave_translator:uav_writedata
	signal capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address                    : std_logic_vector(28 downto 0);  -- capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_address -> capt3_0_avalon_parallel_port_slave_translator:uav_address
	signal capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write                      : std_logic;                      -- capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_write -> capt3_0_avalon_parallel_port_slave_translator:uav_write
	signal capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock                       : std_logic;                      -- capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_lock -> capt3_0_avalon_parallel_port_slave_translator:uav_lock
	signal capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read                       : std_logic;                      -- capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_read -> capt3_0_avalon_parallel_port_slave_translator:uav_read
	signal capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata                   : std_logic_vector(31 downto 0);  -- capt3_0_avalon_parallel_port_slave_translator:uav_readdata -> capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid              : std_logic;                      -- capt3_0_avalon_parallel_port_slave_translator:uav_readdatavalid -> capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess                : std_logic;                      -- capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> capt3_0_avalon_parallel_port_slave_translator:uav_debugaccess
	signal capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable                 : std_logic_vector(3 downto 0);   -- capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> capt3_0_avalon_parallel_port_slave_translator:uav_byteenable
	signal capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket         : std_logic;                      -- capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid               : std_logic;                      -- capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket       : std_logic;                      -- capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data                : std_logic_vector(102 downto 0); -- capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready               : std_logic;                      -- capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket      : std_logic;                      -- capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid            : std_logic;                      -- capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket    : std_logic;                      -- capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data             : std_logic_vector(102 downto 0); -- capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready            : std_logic;                      -- capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid          : std_logic;                      -- capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data           : std_logic_vector(33 downto 0);  -- capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready          : std_logic;                      -- capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest                : std_logic;                      -- capt6_4_avalon_parallel_port_slave_translator:uav_waitrequest -> capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount                 : std_logic_vector(2 downto 0);   -- capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> capt6_4_avalon_parallel_port_slave_translator:uav_burstcount
	signal capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata                  : std_logic_vector(31 downto 0);  -- capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> capt6_4_avalon_parallel_port_slave_translator:uav_writedata
	signal capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address                    : std_logic_vector(28 downto 0);  -- capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_address -> capt6_4_avalon_parallel_port_slave_translator:uav_address
	signal capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write                      : std_logic;                      -- capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_write -> capt6_4_avalon_parallel_port_slave_translator:uav_write
	signal capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock                       : std_logic;                      -- capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_lock -> capt6_4_avalon_parallel_port_slave_translator:uav_lock
	signal capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read                       : std_logic;                      -- capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_read -> capt6_4_avalon_parallel_port_slave_translator:uav_read
	signal capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata                   : std_logic_vector(31 downto 0);  -- capt6_4_avalon_parallel_port_slave_translator:uav_readdata -> capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid              : std_logic;                      -- capt6_4_avalon_parallel_port_slave_translator:uav_readdatavalid -> capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess                : std_logic;                      -- capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> capt6_4_avalon_parallel_port_slave_translator:uav_debugaccess
	signal capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable                 : std_logic_vector(3 downto 0);   -- capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> capt6_4_avalon_parallel_port_slave_translator:uav_byteenable
	signal capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket         : std_logic;                      -- capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid               : std_logic;                      -- capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket       : std_logic;                      -- capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data                : std_logic_vector(102 downto 0); -- capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready               : std_logic;                      -- capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket      : std_logic;                      -- capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid            : std_logic;                      -- capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket    : std_logic;                      -- capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data             : std_logic_vector(102 downto 0); -- capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready            : std_logic;                      -- capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid          : std_logic;                      -- capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data           : std_logic_vector(33 downto 0);  -- capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready          : std_logic;                      -- capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket                           : std_logic;                      -- CPU_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	signal cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid                                 : std_logic;                      -- CPU_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	signal cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket                         : std_logic;                      -- CPU_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	signal cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data                                  : std_logic_vector(101 downto 0); -- CPU_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	signal cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready                                 : std_logic;                      -- addr_router:sink_ready -> CPU_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	signal cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket                                  : std_logic;                      -- CPU_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	signal cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid                                        : std_logic;                      -- CPU_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	signal cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket                                : std_logic;                      -- CPU_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	signal cpu_data_master_translator_avalon_universal_master_0_agent_cp_data                                         : std_logic_vector(101 downto 0); -- CPU_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	signal cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready                                        : std_logic;                      -- addr_router_001:sink_ready -> CPU_data_master_translator_avalon_universal_master_0_agent:cp_ready
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket                             : std_logic;                      -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid                                   : std_logic;                      -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket                           : std_logic;                      -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data                                    : std_logic_vector(101 downto 0); -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready                                   : std_logic;                      -- id_router:sink_ready -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                          : std_logic;                      -- SDRAM_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid                                                : std_logic;                      -- SDRAM_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                        : std_logic;                      -- SDRAM_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rp_data                                                 : std_logic_vector(83 downto 0);  -- SDRAM_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready                                                : std_logic;                      -- id_router_001:sink_ready -> SDRAM_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                 : std_logic;                      -- Interval_timer_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	signal interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid                                       : std_logic;                      -- Interval_timer_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	signal interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                               : std_logic;                      -- Interval_timer_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	signal interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_data                                        : std_logic_vector(101 downto 0); -- Interval_timer_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	signal interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready                                       : std_logic;                      -- id_router_002:sink_ready -> Interval_timer_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket                               : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid                                     : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket                             : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data                                      : std_logic_vector(101 downto 0); -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready                                     : std_logic;                      -- id_router_003:sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket                       : std_logic;                      -- JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid                             : std_logic;                      -- JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket                     : std_logic;                      -- JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data                              : std_logic_vector(101 downto 0); -- JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready                             : std_logic;                      -- id_router_004:sink_ready -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket             : std_logic;                      -- CTR_MOTEUR_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	signal ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid                   : std_logic;                      -- CTR_MOTEUR_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	signal ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket           : std_logic;                      -- CTR_MOTEUR_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	signal ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data                    : std_logic_vector(101 downto 0); -- CTR_MOTEUR_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	signal ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready                   : std_logic;                      -- id_router_005:sink_ready -> CTR_MOTEUR_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket                : std_logic;                      -- capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	signal capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid                      : std_logic;                      -- capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	signal capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket              : std_logic;                      -- capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	signal capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data                       : std_logic_vector(101 downto 0); -- capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	signal capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready                      : std_logic;                      -- id_router_006:sink_ready -> capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket                : std_logic;                      -- capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	signal capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid                      : std_logic;                      -- capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	signal capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket              : std_logic;                      -- capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	signal capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data                       : std_logic_vector(101 downto 0); -- capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	signal capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready                      : std_logic;                      -- id_router_007:sink_ready -> capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal addr_router_src_endofpacket                                                                                : std_logic;                      -- addr_router:src_endofpacket -> limiter:cmd_sink_endofpacket
	signal addr_router_src_valid                                                                                      : std_logic;                      -- addr_router:src_valid -> limiter:cmd_sink_valid
	signal addr_router_src_startofpacket                                                                              : std_logic;                      -- addr_router:src_startofpacket -> limiter:cmd_sink_startofpacket
	signal addr_router_src_data                                                                                       : std_logic_vector(101 downto 0); -- addr_router:src_data -> limiter:cmd_sink_data
	signal addr_router_src_channel                                                                                    : std_logic_vector(7 downto 0);   -- addr_router:src_channel -> limiter:cmd_sink_channel
	signal addr_router_src_ready                                                                                      : std_logic;                      -- limiter:cmd_sink_ready -> addr_router:src_ready
	signal limiter_rsp_src_endofpacket                                                                                : std_logic;                      -- limiter:rsp_src_endofpacket -> CPU_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal limiter_rsp_src_valid                                                                                      : std_logic;                      -- limiter:rsp_src_valid -> CPU_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	signal limiter_rsp_src_startofpacket                                                                              : std_logic;                      -- limiter:rsp_src_startofpacket -> CPU_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal limiter_rsp_src_data                                                                                       : std_logic_vector(101 downto 0); -- limiter:rsp_src_data -> CPU_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	signal limiter_rsp_src_channel                                                                                    : std_logic_vector(7 downto 0);   -- limiter:rsp_src_channel -> CPU_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	signal limiter_rsp_src_ready                                                                                      : std_logic;                      -- CPU_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	signal burst_adapter_source0_endofpacket                                                                          : std_logic;                      -- burst_adapter:source0_endofpacket -> SDRAM_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal burst_adapter_source0_valid                                                                                : std_logic;                      -- burst_adapter:source0_valid -> SDRAM_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal burst_adapter_source0_startofpacket                                                                        : std_logic;                      -- burst_adapter:source0_startofpacket -> SDRAM_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal burst_adapter_source0_data                                                                                 : std_logic_vector(83 downto 0);  -- burst_adapter:source0_data -> SDRAM_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal burst_adapter_source0_ready                                                                                : std_logic;                      -- SDRAM_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	signal burst_adapter_source0_channel                                                                              : std_logic_vector(7 downto 0);   -- burst_adapter:source0_channel -> SDRAM_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal rst_controller_reset_out_reset                                                                             : std_logic;                      -- rst_controller:reset_out -> [CPU_data_master_translator:reset, CPU_data_master_translator_avalon_universal_master_0_agent:reset, CPU_instruction_master_translator:reset, CPU_instruction_master_translator_avalon_universal_master_0_agent:reset, CPU_jtag_debug_module_translator:reset, CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Interval_timer_s1_translator:reset, Interval_timer_s1_translator_avalon_universal_slave_0_agent:reset, Interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, JTAG_UART_avalon_jtag_slave_translator:reset, JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, SDRAM_s1_translator:reset, SDRAM_s1_translator_avalon_universal_slave_0_agent:reset, SDRAM_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, SDRAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, addr_router:reset, addr_router_001:reset, burst_adapter:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, irq_mapper:reset, limiter:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, rst_controller_reset_out_reset:in, sysid_control_slave_translator:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, width_adapter:reset, width_adapter_001:reset]
	signal rst_controller_001_reset_out_reset                                                                         : std_logic;                      -- rst_controller_001:reset_out -> External_Clocks:reset
	signal cmd_xbar_demux_src0_endofpacket                                                                            : std_logic;                      -- cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	signal cmd_xbar_demux_src0_valid                                                                                  : std_logic;                      -- cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	signal cmd_xbar_demux_src0_startofpacket                                                                          : std_logic;                      -- cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	signal cmd_xbar_demux_src0_data                                                                                   : std_logic_vector(101 downto 0); -- cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	signal cmd_xbar_demux_src0_channel                                                                                : std_logic_vector(7 downto 0);   -- cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	signal cmd_xbar_demux_src0_ready                                                                                  : std_logic;                      -- cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	signal cmd_xbar_demux_src1_endofpacket                                                                            : std_logic;                      -- cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	signal cmd_xbar_demux_src1_valid                                                                                  : std_logic;                      -- cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	signal cmd_xbar_demux_src1_startofpacket                                                                          : std_logic;                      -- cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	signal cmd_xbar_demux_src1_data                                                                                   : std_logic_vector(101 downto 0); -- cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	signal cmd_xbar_demux_src1_channel                                                                                : std_logic_vector(7 downto 0);   -- cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	signal cmd_xbar_demux_src1_ready                                                                                  : std_logic;                      -- cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	signal cmd_xbar_demux_001_src0_endofpacket                                                                        : std_logic;                      -- cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	signal cmd_xbar_demux_001_src0_valid                                                                              : std_logic;                      -- cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	signal cmd_xbar_demux_001_src0_startofpacket                                                                      : std_logic;                      -- cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	signal cmd_xbar_demux_001_src0_data                                                                               : std_logic_vector(101 downto 0); -- cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	signal cmd_xbar_demux_001_src0_channel                                                                            : std_logic_vector(7 downto 0);   -- cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	signal cmd_xbar_demux_001_src0_ready                                                                              : std_logic;                      -- cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	signal cmd_xbar_demux_001_src1_endofpacket                                                                        : std_logic;                      -- cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	signal cmd_xbar_demux_001_src1_valid                                                                              : std_logic;                      -- cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	signal cmd_xbar_demux_001_src1_startofpacket                                                                      : std_logic;                      -- cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	signal cmd_xbar_demux_001_src1_data                                                                               : std_logic_vector(101 downto 0); -- cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	signal cmd_xbar_demux_001_src1_channel                                                                            : std_logic_vector(7 downto 0);   -- cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	signal cmd_xbar_demux_001_src1_ready                                                                              : std_logic;                      -- cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	signal cmd_xbar_demux_001_src2_endofpacket                                                                        : std_logic;                      -- cmd_xbar_demux_001:src2_endofpacket -> Interval_timer_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src2_valid                                                                              : std_logic;                      -- cmd_xbar_demux_001:src2_valid -> Interval_timer_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src2_startofpacket                                                                      : std_logic;                      -- cmd_xbar_demux_001:src2_startofpacket -> Interval_timer_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src2_data                                                                               : std_logic_vector(101 downto 0); -- cmd_xbar_demux_001:src2_data -> Interval_timer_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src2_channel                                                                            : std_logic_vector(7 downto 0);   -- cmd_xbar_demux_001:src2_channel -> Interval_timer_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src3_endofpacket                                                                        : std_logic;                      -- cmd_xbar_demux_001:src3_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src3_valid                                                                              : std_logic;                      -- cmd_xbar_demux_001:src3_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src3_startofpacket                                                                      : std_logic;                      -- cmd_xbar_demux_001:src3_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src3_data                                                                               : std_logic_vector(101 downto 0); -- cmd_xbar_demux_001:src3_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src3_channel                                                                            : std_logic_vector(7 downto 0);   -- cmd_xbar_demux_001:src3_channel -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src4_endofpacket                                                                        : std_logic;                      -- cmd_xbar_demux_001:src4_endofpacket -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src4_valid                                                                              : std_logic;                      -- cmd_xbar_demux_001:src4_valid -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src4_startofpacket                                                                      : std_logic;                      -- cmd_xbar_demux_001:src4_startofpacket -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src4_data                                                                               : std_logic_vector(101 downto 0); -- cmd_xbar_demux_001:src4_data -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src4_channel                                                                            : std_logic_vector(7 downto 0);   -- cmd_xbar_demux_001:src4_channel -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src5_endofpacket                                                                        : std_logic;                      -- cmd_xbar_demux_001:src5_endofpacket -> CTR_MOTEUR_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src5_valid                                                                              : std_logic;                      -- cmd_xbar_demux_001:src5_valid -> CTR_MOTEUR_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src5_startofpacket                                                                      : std_logic;                      -- cmd_xbar_demux_001:src5_startofpacket -> CTR_MOTEUR_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src5_data                                                                               : std_logic_vector(101 downto 0); -- cmd_xbar_demux_001:src5_data -> CTR_MOTEUR_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src5_channel                                                                            : std_logic_vector(7 downto 0);   -- cmd_xbar_demux_001:src5_channel -> CTR_MOTEUR_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src6_endofpacket                                                                        : std_logic;                      -- cmd_xbar_demux_001:src6_endofpacket -> capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src6_valid                                                                              : std_logic;                      -- cmd_xbar_demux_001:src6_valid -> capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src6_startofpacket                                                                      : std_logic;                      -- cmd_xbar_demux_001:src6_startofpacket -> capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src6_data                                                                               : std_logic_vector(101 downto 0); -- cmd_xbar_demux_001:src6_data -> capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src6_channel                                                                            : std_logic_vector(7 downto 0);   -- cmd_xbar_demux_001:src6_channel -> capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src7_endofpacket                                                                        : std_logic;                      -- cmd_xbar_demux_001:src7_endofpacket -> capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src7_valid                                                                              : std_logic;                      -- cmd_xbar_demux_001:src7_valid -> capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src7_startofpacket                                                                      : std_logic;                      -- cmd_xbar_demux_001:src7_startofpacket -> capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src7_data                                                                               : std_logic_vector(101 downto 0); -- cmd_xbar_demux_001:src7_data -> capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src7_channel                                                                            : std_logic_vector(7 downto 0);   -- cmd_xbar_demux_001:src7_channel -> capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal rsp_xbar_demux_src0_endofpacket                                                                            : std_logic;                      -- rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	signal rsp_xbar_demux_src0_valid                                                                                  : std_logic;                      -- rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	signal rsp_xbar_demux_src0_startofpacket                                                                          : std_logic;                      -- rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	signal rsp_xbar_demux_src0_data                                                                                   : std_logic_vector(101 downto 0); -- rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	signal rsp_xbar_demux_src0_channel                                                                                : std_logic_vector(7 downto 0);   -- rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	signal rsp_xbar_demux_src0_ready                                                                                  : std_logic;                      -- rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	signal rsp_xbar_demux_src1_endofpacket                                                                            : std_logic;                      -- rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	signal rsp_xbar_demux_src1_valid                                                                                  : std_logic;                      -- rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	signal rsp_xbar_demux_src1_startofpacket                                                                          : std_logic;                      -- rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	signal rsp_xbar_demux_src1_data                                                                                   : std_logic_vector(101 downto 0); -- rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	signal rsp_xbar_demux_src1_channel                                                                                : std_logic_vector(7 downto 0);   -- rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	signal rsp_xbar_demux_src1_ready                                                                                  : std_logic;                      -- rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	signal rsp_xbar_demux_001_src0_endofpacket                                                                        : std_logic;                      -- rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	signal rsp_xbar_demux_001_src0_valid                                                                              : std_logic;                      -- rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	signal rsp_xbar_demux_001_src0_startofpacket                                                                      : std_logic;                      -- rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	signal rsp_xbar_demux_001_src0_data                                                                               : std_logic_vector(101 downto 0); -- rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	signal rsp_xbar_demux_001_src0_channel                                                                            : std_logic_vector(7 downto 0);   -- rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	signal rsp_xbar_demux_001_src0_ready                                                                              : std_logic;                      -- rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	signal rsp_xbar_demux_001_src1_endofpacket                                                                        : std_logic;                      -- rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	signal rsp_xbar_demux_001_src1_valid                                                                              : std_logic;                      -- rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	signal rsp_xbar_demux_001_src1_startofpacket                                                                      : std_logic;                      -- rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	signal rsp_xbar_demux_001_src1_data                                                                               : std_logic_vector(101 downto 0); -- rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	signal rsp_xbar_demux_001_src1_channel                                                                            : std_logic_vector(7 downto 0);   -- rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	signal rsp_xbar_demux_001_src1_ready                                                                              : std_logic;                      -- rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	signal rsp_xbar_demux_002_src0_endofpacket                                                                        : std_logic;                      -- rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	signal rsp_xbar_demux_002_src0_valid                                                                              : std_logic;                      -- rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux_001:sink2_valid
	signal rsp_xbar_demux_002_src0_startofpacket                                                                      : std_logic;                      -- rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	signal rsp_xbar_demux_002_src0_data                                                                               : std_logic_vector(101 downto 0); -- rsp_xbar_demux_002:src0_data -> rsp_xbar_mux_001:sink2_data
	signal rsp_xbar_demux_002_src0_channel                                                                            : std_logic_vector(7 downto 0);   -- rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux_001:sink2_channel
	signal rsp_xbar_demux_002_src0_ready                                                                              : std_logic;                      -- rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_002:src0_ready
	signal rsp_xbar_demux_003_src0_endofpacket                                                                        : std_logic;                      -- rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	signal rsp_xbar_demux_003_src0_valid                                                                              : std_logic;                      -- rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux_001:sink3_valid
	signal rsp_xbar_demux_003_src0_startofpacket                                                                      : std_logic;                      -- rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	signal rsp_xbar_demux_003_src0_data                                                                               : std_logic_vector(101 downto 0); -- rsp_xbar_demux_003:src0_data -> rsp_xbar_mux_001:sink3_data
	signal rsp_xbar_demux_003_src0_channel                                                                            : std_logic_vector(7 downto 0);   -- rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux_001:sink3_channel
	signal rsp_xbar_demux_003_src0_ready                                                                              : std_logic;                      -- rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_003:src0_ready
	signal rsp_xbar_demux_004_src0_endofpacket                                                                        : std_logic;                      -- rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	signal rsp_xbar_demux_004_src0_valid                                                                              : std_logic;                      -- rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux_001:sink4_valid
	signal rsp_xbar_demux_004_src0_startofpacket                                                                      : std_logic;                      -- rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	signal rsp_xbar_demux_004_src0_data                                                                               : std_logic_vector(101 downto 0); -- rsp_xbar_demux_004:src0_data -> rsp_xbar_mux_001:sink4_data
	signal rsp_xbar_demux_004_src0_channel                                                                            : std_logic_vector(7 downto 0);   -- rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux_001:sink4_channel
	signal rsp_xbar_demux_004_src0_ready                                                                              : std_logic;                      -- rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_004:src0_ready
	signal rsp_xbar_demux_005_src0_endofpacket                                                                        : std_logic;                      -- rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	signal rsp_xbar_demux_005_src0_valid                                                                              : std_logic;                      -- rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux_001:sink5_valid
	signal rsp_xbar_demux_005_src0_startofpacket                                                                      : std_logic;                      -- rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	signal rsp_xbar_demux_005_src0_data                                                                               : std_logic_vector(101 downto 0); -- rsp_xbar_demux_005:src0_data -> rsp_xbar_mux_001:sink5_data
	signal rsp_xbar_demux_005_src0_channel                                                                            : std_logic_vector(7 downto 0);   -- rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux_001:sink5_channel
	signal rsp_xbar_demux_005_src0_ready                                                                              : std_logic;                      -- rsp_xbar_mux_001:sink5_ready -> rsp_xbar_demux_005:src0_ready
	signal rsp_xbar_demux_006_src0_endofpacket                                                                        : std_logic;                      -- rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux_001:sink6_endofpacket
	signal rsp_xbar_demux_006_src0_valid                                                                              : std_logic;                      -- rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux_001:sink6_valid
	signal rsp_xbar_demux_006_src0_startofpacket                                                                      : std_logic;                      -- rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux_001:sink6_startofpacket
	signal rsp_xbar_demux_006_src0_data                                                                               : std_logic_vector(101 downto 0); -- rsp_xbar_demux_006:src0_data -> rsp_xbar_mux_001:sink6_data
	signal rsp_xbar_demux_006_src0_channel                                                                            : std_logic_vector(7 downto 0);   -- rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux_001:sink6_channel
	signal rsp_xbar_demux_006_src0_ready                                                                              : std_logic;                      -- rsp_xbar_mux_001:sink6_ready -> rsp_xbar_demux_006:src0_ready
	signal rsp_xbar_demux_007_src0_endofpacket                                                                        : std_logic;                      -- rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux_001:sink7_endofpacket
	signal rsp_xbar_demux_007_src0_valid                                                                              : std_logic;                      -- rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux_001:sink7_valid
	signal rsp_xbar_demux_007_src0_startofpacket                                                                      : std_logic;                      -- rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux_001:sink7_startofpacket
	signal rsp_xbar_demux_007_src0_data                                                                               : std_logic_vector(101 downto 0); -- rsp_xbar_demux_007:src0_data -> rsp_xbar_mux_001:sink7_data
	signal rsp_xbar_demux_007_src0_channel                                                                            : std_logic_vector(7 downto 0);   -- rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux_001:sink7_channel
	signal rsp_xbar_demux_007_src0_ready                                                                              : std_logic;                      -- rsp_xbar_mux_001:sink7_ready -> rsp_xbar_demux_007:src0_ready
	signal limiter_cmd_src_endofpacket                                                                                : std_logic;                      -- limiter:cmd_src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	signal limiter_cmd_src_startofpacket                                                                              : std_logic;                      -- limiter:cmd_src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	signal limiter_cmd_src_data                                                                                       : std_logic_vector(101 downto 0); -- limiter:cmd_src_data -> cmd_xbar_demux:sink_data
	signal limiter_cmd_src_channel                                                                                    : std_logic_vector(7 downto 0);   -- limiter:cmd_src_channel -> cmd_xbar_demux:sink_channel
	signal limiter_cmd_src_ready                                                                                      : std_logic;                      -- cmd_xbar_demux:sink_ready -> limiter:cmd_src_ready
	signal rsp_xbar_mux_src_endofpacket                                                                               : std_logic;                      -- rsp_xbar_mux:src_endofpacket -> limiter:rsp_sink_endofpacket
	signal rsp_xbar_mux_src_valid                                                                                     : std_logic;                      -- rsp_xbar_mux:src_valid -> limiter:rsp_sink_valid
	signal rsp_xbar_mux_src_startofpacket                                                                             : std_logic;                      -- rsp_xbar_mux:src_startofpacket -> limiter:rsp_sink_startofpacket
	signal rsp_xbar_mux_src_data                                                                                      : std_logic_vector(101 downto 0); -- rsp_xbar_mux:src_data -> limiter:rsp_sink_data
	signal rsp_xbar_mux_src_channel                                                                                   : std_logic_vector(7 downto 0);   -- rsp_xbar_mux:src_channel -> limiter:rsp_sink_channel
	signal rsp_xbar_mux_src_ready                                                                                     : std_logic;                      -- limiter:rsp_sink_ready -> rsp_xbar_mux:src_ready
	signal addr_router_001_src_endofpacket                                                                            : std_logic;                      -- addr_router_001:src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	signal addr_router_001_src_valid                                                                                  : std_logic;                      -- addr_router_001:src_valid -> cmd_xbar_demux_001:sink_valid
	signal addr_router_001_src_startofpacket                                                                          : std_logic;                      -- addr_router_001:src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	signal addr_router_001_src_data                                                                                   : std_logic_vector(101 downto 0); -- addr_router_001:src_data -> cmd_xbar_demux_001:sink_data
	signal addr_router_001_src_channel                                                                                : std_logic_vector(7 downto 0);   -- addr_router_001:src_channel -> cmd_xbar_demux_001:sink_channel
	signal addr_router_001_src_ready                                                                                  : std_logic;                      -- cmd_xbar_demux_001:sink_ready -> addr_router_001:src_ready
	signal rsp_xbar_mux_001_src_endofpacket                                                                           : std_logic;                      -- rsp_xbar_mux_001:src_endofpacket -> CPU_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal rsp_xbar_mux_001_src_valid                                                                                 : std_logic;                      -- rsp_xbar_mux_001:src_valid -> CPU_data_master_translator_avalon_universal_master_0_agent:rp_valid
	signal rsp_xbar_mux_001_src_startofpacket                                                                         : std_logic;                      -- rsp_xbar_mux_001:src_startofpacket -> CPU_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal rsp_xbar_mux_001_src_data                                                                                  : std_logic_vector(101 downto 0); -- rsp_xbar_mux_001:src_data -> CPU_data_master_translator_avalon_universal_master_0_agent:rp_data
	signal rsp_xbar_mux_001_src_channel                                                                               : std_logic_vector(7 downto 0);   -- rsp_xbar_mux_001:src_channel -> CPU_data_master_translator_avalon_universal_master_0_agent:rp_channel
	signal rsp_xbar_mux_001_src_ready                                                                                 : std_logic;                      -- CPU_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_001:src_ready
	signal cmd_xbar_mux_src_endofpacket                                                                               : std_logic;                      -- cmd_xbar_mux:src_endofpacket -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_src_valid                                                                                     : std_logic;                      -- cmd_xbar_mux:src_valid -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_src_startofpacket                                                                             : std_logic;                      -- cmd_xbar_mux:src_startofpacket -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_src_data                                                                                      : std_logic_vector(101 downto 0); -- cmd_xbar_mux:src_data -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_src_channel                                                                                   : std_logic_vector(7 downto 0);   -- cmd_xbar_mux:src_channel -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_src_ready                                                                                     : std_logic;                      -- CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	signal id_router_src_endofpacket                                                                                  : std_logic;                      -- id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	signal id_router_src_valid                                                                                        : std_logic;                      -- id_router:src_valid -> rsp_xbar_demux:sink_valid
	signal id_router_src_startofpacket                                                                                : std_logic;                      -- id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	signal id_router_src_data                                                                                         : std_logic_vector(101 downto 0); -- id_router:src_data -> rsp_xbar_demux:sink_data
	signal id_router_src_channel                                                                                      : std_logic_vector(7 downto 0);   -- id_router:src_channel -> rsp_xbar_demux:sink_channel
	signal id_router_src_ready                                                                                        : std_logic;                      -- rsp_xbar_demux:sink_ready -> id_router:src_ready
	signal cmd_xbar_demux_001_src2_ready                                                                              : std_logic;                      -- Interval_timer_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src2_ready
	signal id_router_002_src_endofpacket                                                                              : std_logic;                      -- id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	signal id_router_002_src_valid                                                                                    : std_logic;                      -- id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	signal id_router_002_src_startofpacket                                                                            : std_logic;                      -- id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	signal id_router_002_src_data                                                                                     : std_logic_vector(101 downto 0); -- id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	signal id_router_002_src_channel                                                                                  : std_logic_vector(7 downto 0);   -- id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	signal id_router_002_src_ready                                                                                    : std_logic;                      -- rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	signal cmd_xbar_demux_001_src3_ready                                                                              : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src3_ready
	signal id_router_003_src_endofpacket                                                                              : std_logic;                      -- id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	signal id_router_003_src_valid                                                                                    : std_logic;                      -- id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	signal id_router_003_src_startofpacket                                                                            : std_logic;                      -- id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	signal id_router_003_src_data                                                                                     : std_logic_vector(101 downto 0); -- id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	signal id_router_003_src_channel                                                                                  : std_logic_vector(7 downto 0);   -- id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	signal id_router_003_src_ready                                                                                    : std_logic;                      -- rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	signal cmd_xbar_demux_001_src4_ready                                                                              : std_logic;                      -- JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src4_ready
	signal id_router_004_src_endofpacket                                                                              : std_logic;                      -- id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	signal id_router_004_src_valid                                                                                    : std_logic;                      -- id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	signal id_router_004_src_startofpacket                                                                            : std_logic;                      -- id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	signal id_router_004_src_data                                                                                     : std_logic_vector(101 downto 0); -- id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	signal id_router_004_src_channel                                                                                  : std_logic_vector(7 downto 0);   -- id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	signal id_router_004_src_ready                                                                                    : std_logic;                      -- rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	signal cmd_xbar_demux_001_src5_ready                                                                              : std_logic;                      -- CTR_MOTEUR_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src5_ready
	signal id_router_005_src_endofpacket                                                                              : std_logic;                      -- id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	signal id_router_005_src_valid                                                                                    : std_logic;                      -- id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	signal id_router_005_src_startofpacket                                                                            : std_logic;                      -- id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	signal id_router_005_src_data                                                                                     : std_logic_vector(101 downto 0); -- id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	signal id_router_005_src_channel                                                                                  : std_logic_vector(7 downto 0);   -- id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	signal id_router_005_src_ready                                                                                    : std_logic;                      -- rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	signal cmd_xbar_demux_001_src6_ready                                                                              : std_logic;                      -- capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src6_ready
	signal id_router_006_src_endofpacket                                                                              : std_logic;                      -- id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	signal id_router_006_src_valid                                                                                    : std_logic;                      -- id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	signal id_router_006_src_startofpacket                                                                            : std_logic;                      -- id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	signal id_router_006_src_data                                                                                     : std_logic_vector(101 downto 0); -- id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	signal id_router_006_src_channel                                                                                  : std_logic_vector(7 downto 0);   -- id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	signal id_router_006_src_ready                                                                                    : std_logic;                      -- rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	signal cmd_xbar_demux_001_src7_ready                                                                              : std_logic;                      -- capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src7_ready
	signal id_router_007_src_endofpacket                                                                              : std_logic;                      -- id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	signal id_router_007_src_valid                                                                                    : std_logic;                      -- id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	signal id_router_007_src_startofpacket                                                                            : std_logic;                      -- id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	signal id_router_007_src_data                                                                                     : std_logic_vector(101 downto 0); -- id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	signal id_router_007_src_channel                                                                                  : std_logic_vector(7 downto 0);   -- id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	signal id_router_007_src_ready                                                                                    : std_logic;                      -- rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	signal cmd_xbar_mux_001_src_endofpacket                                                                           : std_logic;                      -- cmd_xbar_mux_001:src_endofpacket -> width_adapter:in_endofpacket
	signal cmd_xbar_mux_001_src_valid                                                                                 : std_logic;                      -- cmd_xbar_mux_001:src_valid -> width_adapter:in_valid
	signal cmd_xbar_mux_001_src_startofpacket                                                                         : std_logic;                      -- cmd_xbar_mux_001:src_startofpacket -> width_adapter:in_startofpacket
	signal cmd_xbar_mux_001_src_data                                                                                  : std_logic_vector(101 downto 0); -- cmd_xbar_mux_001:src_data -> width_adapter:in_data
	signal cmd_xbar_mux_001_src_channel                                                                               : std_logic_vector(7 downto 0);   -- cmd_xbar_mux_001:src_channel -> width_adapter:in_channel
	signal cmd_xbar_mux_001_src_ready                                                                                 : std_logic;                      -- width_adapter:in_ready -> cmd_xbar_mux_001:src_ready
	signal width_adapter_src_endofpacket                                                                              : std_logic;                      -- width_adapter:out_endofpacket -> burst_adapter:sink0_endofpacket
	signal width_adapter_src_valid                                                                                    : std_logic;                      -- width_adapter:out_valid -> burst_adapter:sink0_valid
	signal width_adapter_src_startofpacket                                                                            : std_logic;                      -- width_adapter:out_startofpacket -> burst_adapter:sink0_startofpacket
	signal width_adapter_src_data                                                                                     : std_logic_vector(83 downto 0);  -- width_adapter:out_data -> burst_adapter:sink0_data
	signal width_adapter_src_ready                                                                                    : std_logic;                      -- burst_adapter:sink0_ready -> width_adapter:out_ready
	signal width_adapter_src_channel                                                                                  : std_logic_vector(7 downto 0);   -- width_adapter:out_channel -> burst_adapter:sink0_channel
	signal id_router_001_src_endofpacket                                                                              : std_logic;                      -- id_router_001:src_endofpacket -> width_adapter_001:in_endofpacket
	signal id_router_001_src_valid                                                                                    : std_logic;                      -- id_router_001:src_valid -> width_adapter_001:in_valid
	signal id_router_001_src_startofpacket                                                                            : std_logic;                      -- id_router_001:src_startofpacket -> width_adapter_001:in_startofpacket
	signal id_router_001_src_data                                                                                     : std_logic_vector(83 downto 0);  -- id_router_001:src_data -> width_adapter_001:in_data
	signal id_router_001_src_channel                                                                                  : std_logic_vector(7 downto 0);   -- id_router_001:src_channel -> width_adapter_001:in_channel
	signal id_router_001_src_ready                                                                                    : std_logic;                      -- width_adapter_001:in_ready -> id_router_001:src_ready
	signal width_adapter_001_src_endofpacket                                                                          : std_logic;                      -- width_adapter_001:out_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	signal width_adapter_001_src_valid                                                                                : std_logic;                      -- width_adapter_001:out_valid -> rsp_xbar_demux_001:sink_valid
	signal width_adapter_001_src_startofpacket                                                                        : std_logic;                      -- width_adapter_001:out_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	signal width_adapter_001_src_data                                                                                 : std_logic_vector(101 downto 0); -- width_adapter_001:out_data -> rsp_xbar_demux_001:sink_data
	signal width_adapter_001_src_ready                                                                                : std_logic;                      -- rsp_xbar_demux_001:sink_ready -> width_adapter_001:out_ready
	signal width_adapter_001_src_channel                                                                              : std_logic_vector(7 downto 0);   -- width_adapter_001:out_channel -> rsp_xbar_demux_001:sink_channel
	signal limiter_cmd_valid_data                                                                                     : std_logic_vector(7 downto 0);   -- limiter:cmd_src_valid -> cmd_xbar_demux:sink_valid
	signal irq_mapper_receiver0_irq                                                                                   : std_logic;                      -- JTAG_UART:av_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                                                                   : std_logic;                      -- Interval_timer:irq -> irq_mapper:receiver1_irq
	signal cpu_d_irq_irq                                                                                              : std_logic_vector(31 downto 0);  -- irq_mapper:sender_irq -> CPU:d_irq
	signal reset_n_ports_inv                                                                                          : std_logic;                      -- reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0]
	signal sdram_s1_translator_avalon_anti_slave_0_write_ports_inv                                                    : std_logic;                      -- sdram_s1_translator_avalon_anti_slave_0_write:inv -> SDRAM:az_wr_n
	signal sdram_s1_translator_avalon_anti_slave_0_read_ports_inv                                                     : std_logic;                      -- sdram_s1_translator_avalon_anti_slave_0_read:inv -> SDRAM:az_rd_n
	signal sdram_s1_translator_avalon_anti_slave_0_byteenable_ports_inv                                               : std_logic_vector(1 downto 0);   -- sdram_s1_translator_avalon_anti_slave_0_byteenable:inv -> SDRAM:az_be_n
	signal interval_timer_s1_translator_avalon_anti_slave_0_write_ports_inv                                           : std_logic;                      -- interval_timer_s1_translator_avalon_anti_slave_0_write:inv -> Interval_timer:write_n
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write_ports_inv                                 : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write:inv -> JTAG_UART:av_write_n
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read_ports_inv                                  : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read:inv -> JTAG_UART:av_read_n
	signal rst_controller_reset_out_reset_ports_inv                                                                   : std_logic;                      -- rst_controller_reset_out_reset:inv -> [CPU:reset_n, Interval_timer:reset_n, JTAG_UART:rst_n, SDRAM:reset_n, sysid:reset_n]

begin

	jtag_uart : component nios_system_JTAG_UART
		port map (
			clk            => external_clocks_sys_clk_clk,                                                --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                                   --             reset.reset_n
			av_chipselect  => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address(0),      --                  .address
			av_read_n      => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read_ports_inv,  --                  .read_n
			av_readdata    => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata,        --                  .readdata
			av_write_n     => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write_ports_inv, --                  .write_n
			av_writedata   => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata,       --                  .writedata
			av_waitrequest => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                                    --               irq.irq
		);

	interval_timer : component nios_system_Interval_timer
		port map (
			clk        => external_clocks_sys_clk_clk,                                      --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                         -- reset.reset_n
			address    => interval_timer_s1_translator_avalon_anti_slave_0_address,         --    s1.address
			writedata  => interval_timer_s1_translator_avalon_anti_slave_0_writedata,       --      .writedata
			readdata   => interval_timer_s1_translator_avalon_anti_slave_0_readdata,        --      .readdata
			chipselect => interval_timer_s1_translator_avalon_anti_slave_0_chipselect,      --      .chipselect
			write_n    => interval_timer_s1_translator_avalon_anti_slave_0_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver1_irq                                          --   irq.irq
		);

	sdram : component nios_system_SDRAM
		port map (
			clk            => external_clocks_sys_clk_clk,                                  --   clk.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,                     -- reset.reset_n
			az_addr        => sdram_s1_translator_avalon_anti_slave_0_address,              --    s1.address
			az_be_n        => sdram_s1_translator_avalon_anti_slave_0_byteenable_ports_inv, --      .byteenable_n
			az_cs          => sdram_s1_translator_avalon_anti_slave_0_chipselect,           --      .chipselect
			az_data        => sdram_s1_translator_avalon_anti_slave_0_writedata,            --      .writedata
			az_rd_n        => sdram_s1_translator_avalon_anti_slave_0_read_ports_inv,       --      .read_n
			az_wr_n        => sdram_s1_translator_avalon_anti_slave_0_write_ports_inv,      --      .write_n
			za_data        => sdram_s1_translator_avalon_anti_slave_0_readdata,             --      .readdata
			za_valid       => sdram_s1_translator_avalon_anti_slave_0_readdatavalid,        --      .readdatavalid
			za_waitrequest => sdram_s1_translator_avalon_anti_slave_0_waitrequest,          --      .waitrequest
			zs_addr        => zs_addr_from_the_SDRAM,                                       --  wire.export
			zs_ba          => zs_ba_from_the_SDRAM,                                         --      .export
			zs_cas_n       => zs_cas_n_from_the_SDRAM,                                      --      .export
			zs_cke         => zs_cke_from_the_SDRAM,                                        --      .export
			zs_cs_n        => zs_cs_n_from_the_SDRAM,                                       --      .export
			zs_dq          => zs_dq_to_and_from_the_SDRAM,                                  --      .export
			zs_dqm         => zs_dqm_from_the_SDRAM,                                        --      .export
			zs_ras_n       => zs_ras_n_from_the_SDRAM,                                      --      .export
			zs_we_n        => zs_we_n_from_the_SDRAM                                        --      .export
		);

	cpu : component nios_system_CPU
		port map (
			clk                                   => external_clocks_sys_clk_clk,                                      --                       clk.clk
			reset_n                               => rst_controller_reset_out_reset_ports_inv,                         --                   reset_n.reset_n
			d_address                             => cpu_data_master_address,                                          --               data_master.address
			d_byteenable                          => cpu_data_master_byteenable,                                       --                          .byteenable
			d_read                                => cpu_data_master_read,                                             --                          .read
			d_readdata                            => cpu_data_master_readdata,                                         --                          .readdata
			d_waitrequest                         => cpu_data_master_waitrequest,                                      --                          .waitrequest
			d_write                               => cpu_data_master_write,                                            --                          .write
			d_writedata                           => cpu_data_master_writedata,                                        --                          .writedata
			jtag_debug_module_debugaccess_to_roms => cpu_data_master_debugaccess,                                      --                          .debugaccess
			i_address                             => cpu_instruction_master_address,                                   --        instruction_master.address
			i_read                                => cpu_instruction_master_read,                                      --                          .read
			i_readdata                            => cpu_instruction_master_readdata,                                  --                          .readdata
			i_waitrequest                         => cpu_instruction_master_waitrequest,                               --                          .waitrequest
			i_readdatavalid                       => cpu_instruction_master_readdatavalid,                             --                          .readdatavalid
			d_irq                                 => cpu_d_irq_irq,                                                    --                     d_irq.irq
			jtag_debug_module_resetrequest        => cpu_jtag_debug_module_reset_reset,                                --   jtag_debug_module_reset.reset
			jtag_debug_module_address             => cpu_jtag_debug_module_translator_avalon_anti_slave_0_address,     --         jtag_debug_module.address
			jtag_debug_module_byteenable          => cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable,  --                          .byteenable
			jtag_debug_module_debugaccess         => cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess, --                          .debugaccess
			jtag_debug_module_read                => cpu_jtag_debug_module_translator_avalon_anti_slave_0_read,        --                          .read
			jtag_debug_module_readdata            => cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata,    --                          .readdata
			jtag_debug_module_waitrequest         => cpu_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest, --                          .waitrequest
			jtag_debug_module_write               => cpu_jtag_debug_module_translator_avalon_anti_slave_0_write,       --                          .write
			jtag_debug_module_writedata           => cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata,   --                          .writedata
			no_ci_readra                          => open                                                              -- custom_instruction_master.readra
		);

	sysid : component nios_system_sysid
		port map (
			clock    => external_clocks_sys_clk_clk,                                   --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,                      --         reset.reset_n
			readdata => sysid_control_slave_translator_avalon_anti_slave_0_readdata,   -- control_slave.readdata
			address  => sysid_control_slave_translator_avalon_anti_slave_0_address(0)  --              .address
		);

	external_clocks : component nios_system_External_Clocks
		port map (
			CLOCK_50    => clk,                                --       clk_in_primary.clk
			reset       => rst_controller_001_reset_out_reset, -- clk_in_primary_reset.reset
			sys_clk     => external_clocks_sys_clk_clk,        --              sys_clk.clk
			sys_reset_n => open,                               --        sys_clk_reset.reset_n
			SDRAM_CLK   => sdram_clk                           --            sdram_clk.clk
		);

	ctr_moteur : component nios_system_CTR_MOTEUR
		port map (
			clk        => external_clocks_sys_clk_clk,                                                     --                clock_reset.clk
			reset      => cpu_jtag_debug_module_reset_reset,                                               --          clock_reset_reset.reset
			address    => ctr_moteur_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address,    -- avalon_parallel_port_slave.address
			byteenable => ctr_moteur_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable, --                           .byteenable
			chipselect => ctr_moteur_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect, --                           .chipselect
			read       => ctr_moteur_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read,       --                           .read
			write      => ctr_moteur_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write,      --                           .write
			writedata  => ctr_moteur_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata,  --                           .writedata
			readdata   => ctr_moteur_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata,   --                           .readdata
			out_port   => omoteurctr_export                                                                --         external_interface.export
		);

	capt3_0 : component nios_system_capt3_0
		port map (
			clk        => external_clocks_sys_clk_clk,                                                  --                clock_reset.clk
			reset      => cpu_jtag_debug_module_reset_reset,                                            --          clock_reset_reset.reset
			address    => capt3_0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address,    -- avalon_parallel_port_slave.address
			byteenable => capt3_0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable, --                           .byteenable
			chipselect => capt3_0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect, --                           .chipselect
			read       => capt3_0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read,       --                           .read
			write      => capt3_0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write,      --                           .write
			writedata  => capt3_0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata,  --                           .writedata
			readdata   => capt3_0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata,   --                           .readdata
			in_port    => capt3_0_signal_export                                                         --         external_interface.export
		);

	capt6_4 : component nios_system_capt3_0
		port map (
			clk        => external_clocks_sys_clk_clk,                                                  --                clock_reset.clk
			reset      => cpu_jtag_debug_module_reset_reset,                                            --          clock_reset_reset.reset
			address    => capt6_4_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address,    -- avalon_parallel_port_slave.address
			byteenable => capt6_4_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable, --                           .byteenable
			chipselect => capt6_4_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect, --                           .chipselect
			read       => capt6_4_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read,       --                           .read
			write      => capt6_4_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write,      --                           .write
			writedata  => capt6_4_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata,  --                           .writedata
			readdata   => capt6_4_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata,   --                           .readdata
			in_port    => capt6_4_signal_export                                                         --         external_interface.export
		);

	cpu_instruction_master_translator : component nios_system_cpu_instruction_master_translator
		generic map (
			AV_ADDRESS_W                => 28,
			AV_DATA_W                   => 32,
			AV_BURSTCOUNT_W             => 1,
			AV_BYTEENABLE_W             => 4,
			UAV_ADDRESS_W               => 29,
			UAV_BURSTCOUNT_W            => 3,
			USE_READ                    => 1,
			USE_WRITE                   => 0,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 0,
			USE_READDATAVALID           => 1,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 4,
			AV_ADDRESS_SYMBOLS          => 1,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 0,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 1,
			AV_REGISTERINCOMINGSIGNALS  => 0
		)
		port map (
			clk                      => external_clocks_sys_clk_clk,                                               --                       clk.clk
			reset                    => rst_controller_reset_out_reset,                                            --                     reset.reset
			uav_address              => cpu_instruction_master_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => cpu_instruction_master_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => cpu_instruction_master_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => cpu_instruction_master_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => cpu_instruction_master_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => cpu_instruction_master_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => cpu_instruction_master_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => cpu_instruction_master_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => cpu_instruction_master_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => cpu_instruction_master_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address               => cpu_instruction_master_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => cpu_instruction_master_waitrequest,                                        --                          .waitrequest
			av_read                  => cpu_instruction_master_read,                                               --                          .read
			av_readdata              => cpu_instruction_master_readdata,                                           --                          .readdata
			av_readdatavalid         => cpu_instruction_master_readdatavalid,                                      --                          .readdatavalid
			av_burstcount            => "1",                                                                       --               (terminated)
			av_byteenable            => "1111",                                                                    --               (terminated)
			av_beginbursttransfer    => '0',                                                                       --               (terminated)
			av_begintransfer         => '0',                                                                       --               (terminated)
			av_chipselect            => '0',                                                                       --               (terminated)
			av_write                 => '0',                                                                       --               (terminated)
			av_writedata             => "00000000000000000000000000000000",                                        --               (terminated)
			av_lock                  => '0',                                                                       --               (terminated)
			av_debugaccess           => '0',                                                                       --               (terminated)
			uav_clken                => open,                                                                      --               (terminated)
			av_clken                 => '1',                                                                       --               (terminated)
			uav_response             => "00",                                                                      --               (terminated)
			av_response              => open,                                                                      --               (terminated)
			uav_writeresponserequest => open,                                                                      --               (terminated)
			uav_writeresponsevalid   => '0',                                                                       --               (terminated)
			av_writeresponserequest  => '0',                                                                       --               (terminated)
			av_writeresponsevalid    => open                                                                       --               (terminated)
		);

	cpu_data_master_translator : component nios_system_cpu_data_master_translator
		generic map (
			AV_ADDRESS_W                => 29,
			AV_DATA_W                   => 32,
			AV_BURSTCOUNT_W             => 1,
			AV_BYTEENABLE_W             => 4,
			UAV_ADDRESS_W               => 29,
			UAV_BURSTCOUNT_W            => 3,
			USE_READ                    => 1,
			USE_WRITE                   => 1,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 0,
			USE_READDATAVALID           => 0,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 4,
			AV_ADDRESS_SYMBOLS          => 1,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 0,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 0,
			AV_REGISTERINCOMINGSIGNALS  => 0
		)
		port map (
			clk                      => external_clocks_sys_clk_clk,                                        --                       clk.clk
			reset                    => rst_controller_reset_out_reset,                                     --                     reset.reset
			uav_address              => cpu_data_master_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => cpu_data_master_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => cpu_data_master_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => cpu_data_master_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => cpu_data_master_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => cpu_data_master_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => cpu_data_master_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => cpu_data_master_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => cpu_data_master_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => cpu_data_master_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => cpu_data_master_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address               => cpu_data_master_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => cpu_data_master_waitrequest,                                        --                          .waitrequest
			av_byteenable            => cpu_data_master_byteenable,                                         --                          .byteenable
			av_read                  => cpu_data_master_read,                                               --                          .read
			av_readdata              => cpu_data_master_readdata,                                           --                          .readdata
			av_write                 => cpu_data_master_write,                                              --                          .write
			av_writedata             => cpu_data_master_writedata,                                          --                          .writedata
			av_debugaccess           => cpu_data_master_debugaccess,                                        --                          .debugaccess
			av_burstcount            => "1",                                                                --               (terminated)
			av_beginbursttransfer    => '0',                                                                --               (terminated)
			av_begintransfer         => '0',                                                                --               (terminated)
			av_chipselect            => '0',                                                                --               (terminated)
			av_readdatavalid         => open,                                                               --               (terminated)
			av_lock                  => '0',                                                                --               (terminated)
			uav_clken                => open,                                                               --               (terminated)
			av_clken                 => '1',                                                                --               (terminated)
			uav_response             => "00",                                                               --               (terminated)
			av_response              => open,                                                               --               (terminated)
			uav_writeresponserequest => open,                                                               --               (terminated)
			uav_writeresponsevalid   => '0',                                                                --               (terminated)
			av_writeresponserequest  => '0',                                                                --               (terminated)
			av_writeresponsevalid    => open                                                                --               (terminated)
		);

	cpu_jtag_debug_module_translator : component nios_system_cpu_jtag_debug_module_translator
		generic map (
			AV_ADDRESS_W                   => 9,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 29,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => external_clocks_sys_clk_clk,                                                      --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                   --                    reset.reset
			uav_address              => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => cpu_jtag_debug_module_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => cpu_jtag_debug_module_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => cpu_jtag_debug_module_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable            => cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_waitrequest           => cpu_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_debugaccess           => cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess,                 --                         .debugaccess
			av_begintransfer         => open,                                                                             --              (terminated)
			av_beginbursttransfer    => open,                                                                             --              (terminated)
			av_burstcount            => open,                                                                             --              (terminated)
			av_readdatavalid         => '0',                                                                              --              (terminated)
			av_writebyteenable       => open,                                                                             --              (terminated)
			av_lock                  => open,                                                                             --              (terminated)
			av_chipselect            => open,                                                                             --              (terminated)
			av_clken                 => open,                                                                             --              (terminated)
			uav_clken                => '0',                                                                              --              (terminated)
			av_outputenable          => open,                                                                             --              (terminated)
			uav_response             => open,                                                                             --              (terminated)
			av_response              => "00",                                                                             --              (terminated)
			uav_writeresponserequest => '0',                                                                              --              (terminated)
			uav_writeresponsevalid   => open,                                                                             --              (terminated)
			av_writeresponserequest  => open,                                                                             --              (terminated)
			av_writeresponsevalid    => '0'                                                                               --              (terminated)
		);

	sdram_s1_translator : component nios_system_sdram_s1_translator
		generic map (
			AV_ADDRESS_W                   => 24,
			AV_DATA_W                      => 16,
			UAV_DATA_W                     => 16,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 2,
			UAV_BYTEENABLE_W               => 2,
			UAV_ADDRESS_W                  => 29,
			UAV_BURSTCOUNT_W               => 2,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 1,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 2,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => external_clocks_sys_clk_clk,                                         --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                      --                    reset.reset
			uav_address              => sdram_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => sdram_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => sdram_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => sdram_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => sdram_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => sdram_s1_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => sdram_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => sdram_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable            => sdram_s1_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_readdatavalid         => sdram_s1_translator_avalon_anti_slave_0_readdatavalid,               --                         .readdatavalid
			av_waitrequest           => sdram_s1_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_chipselect            => sdram_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_begintransfer         => open,                                                                --              (terminated)
			av_beginbursttransfer    => open,                                                                --              (terminated)
			av_burstcount            => open,                                                                --              (terminated)
			av_writebyteenable       => open,                                                                --              (terminated)
			av_lock                  => open,                                                                --              (terminated)
			av_clken                 => open,                                                                --              (terminated)
			uav_clken                => '0',                                                                 --              (terminated)
			av_debugaccess           => open,                                                                --              (terminated)
			av_outputenable          => open,                                                                --              (terminated)
			uav_response             => open,                                                                --              (terminated)
			av_response              => "00",                                                                --              (terminated)
			uav_writeresponserequest => '0',                                                                 --              (terminated)
			uav_writeresponsevalid   => open,                                                                --              (terminated)
			av_writeresponserequest  => open,                                                                --              (terminated)
			av_writeresponsevalid    => '0'                                                                  --              (terminated)
		);

	interval_timer_s1_translator : component nios_system_interval_timer_s1_translator
		generic map (
			AV_ADDRESS_W                   => 3,
			AV_DATA_W                      => 16,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 29,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => external_clocks_sys_clk_clk,                                                  --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                               --                    reset.reset
			uav_address              => interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => interval_timer_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => interval_timer_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => interval_timer_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => interval_timer_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => interval_timer_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                         --              (terminated)
			av_begintransfer         => open,                                                                         --              (terminated)
			av_beginbursttransfer    => open,                                                                         --              (terminated)
			av_burstcount            => open,                                                                         --              (terminated)
			av_byteenable            => open,                                                                         --              (terminated)
			av_readdatavalid         => '0',                                                                          --              (terminated)
			av_waitrequest           => '0',                                                                          --              (terminated)
			av_writebyteenable       => open,                                                                         --              (terminated)
			av_lock                  => open,                                                                         --              (terminated)
			av_clken                 => open,                                                                         --              (terminated)
			uav_clken                => '0',                                                                          --              (terminated)
			av_debugaccess           => open,                                                                         --              (terminated)
			av_outputenable          => open,                                                                         --              (terminated)
			uav_response             => open,                                                                         --              (terminated)
			av_response              => "00",                                                                         --              (terminated)
			uav_writeresponserequest => '0',                                                                          --              (terminated)
			uav_writeresponsevalid   => open,                                                                         --              (terminated)
			av_writeresponserequest  => open,                                                                         --              (terminated)
			av_writeresponsevalid    => '0'                                                                           --              (terminated)
		);

	sysid_control_slave_translator : component nios_system_sysid_control_slave_translator
		generic map (
			AV_ADDRESS_W                   => 1,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 29,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => external_clocks_sys_clk_clk,                                                    --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                 --                    reset.reset
			uav_address              => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => sysid_control_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_readdata              => sysid_control_slave_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_write                 => open,                                                                           --              (terminated)
			av_read                  => open,                                                                           --              (terminated)
			av_writedata             => open,                                                                           --              (terminated)
			av_begintransfer         => open,                                                                           --              (terminated)
			av_beginbursttransfer    => open,                                                                           --              (terminated)
			av_burstcount            => open,                                                                           --              (terminated)
			av_byteenable            => open,                                                                           --              (terminated)
			av_readdatavalid         => '0',                                                                            --              (terminated)
			av_waitrequest           => '0',                                                                            --              (terminated)
			av_writebyteenable       => open,                                                                           --              (terminated)
			av_lock                  => open,                                                                           --              (terminated)
			av_chipselect            => open,                                                                           --              (terminated)
			av_clken                 => open,                                                                           --              (terminated)
			uav_clken                => '0',                                                                            --              (terminated)
			av_debugaccess           => open,                                                                           --              (terminated)
			av_outputenable          => open,                                                                           --              (terminated)
			uav_response             => open,                                                                           --              (terminated)
			av_response              => "00",                                                                           --              (terminated)
			uav_writeresponserequest => '0',                                                                            --              (terminated)
			uav_writeresponsevalid   => open,                                                                           --              (terminated)
			av_writeresponserequest  => open,                                                                           --              (terminated)
			av_writeresponsevalid    => '0'                                                                             --              (terminated)
		);

	jtag_uart_avalon_jtag_slave_translator : component nios_system_jtag_uart_avalon_jtag_slave_translator
		generic map (
			AV_ADDRESS_W                   => 1,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 29,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => external_clocks_sys_clk_clk,                                                            --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                         --                    reset.reset
			uav_address              => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_waitrequest           => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_chipselect            => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_begintransfer         => open,                                                                                   --              (terminated)
			av_beginbursttransfer    => open,                                                                                   --              (terminated)
			av_burstcount            => open,                                                                                   --              (terminated)
			av_byteenable            => open,                                                                                   --              (terminated)
			av_readdatavalid         => '0',                                                                                    --              (terminated)
			av_writebyteenable       => open,                                                                                   --              (terminated)
			av_lock                  => open,                                                                                   --              (terminated)
			av_clken                 => open,                                                                                   --              (terminated)
			uav_clken                => '0',                                                                                    --              (terminated)
			av_debugaccess           => open,                                                                                   --              (terminated)
			av_outputenable          => open,                                                                                   --              (terminated)
			uav_response             => open,                                                                                   --              (terminated)
			av_response              => "00",                                                                                   --              (terminated)
			uav_writeresponserequest => '0',                                                                                    --              (terminated)
			uav_writeresponsevalid   => open,                                                                                   --              (terminated)
			av_writeresponserequest  => open,                                                                                   --              (terminated)
			av_writeresponsevalid    => '0'                                                                                     --              (terminated)
		);

	ctr_moteur_avalon_parallel_port_slave_translator : component nios_system_ctr_moteur_avalon_parallel_port_slave_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 29,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 1,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 0,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => external_clocks_sys_clk_clk,                                                                      --                      clk.clk
			reset                    => cpu_jtag_debug_module_reset_reset,                                                                --                    reset.reset
			uav_address              => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => ctr_moteur_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => ctr_moteur_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => ctr_moteur_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => ctr_moteur_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => ctr_moteur_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable            => ctr_moteur_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_chipselect            => ctr_moteur_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_begintransfer         => open,                                                                                             --              (terminated)
			av_beginbursttransfer    => open,                                                                                             --              (terminated)
			av_burstcount            => open,                                                                                             --              (terminated)
			av_readdatavalid         => '0',                                                                                              --              (terminated)
			av_waitrequest           => '0',                                                                                              --              (terminated)
			av_writebyteenable       => open,                                                                                             --              (terminated)
			av_lock                  => open,                                                                                             --              (terminated)
			av_clken                 => open,                                                                                             --              (terminated)
			uav_clken                => '0',                                                                                              --              (terminated)
			av_debugaccess           => open,                                                                                             --              (terminated)
			av_outputenable          => open,                                                                                             --              (terminated)
			uav_response             => open,                                                                                             --              (terminated)
			av_response              => "00",                                                                                             --              (terminated)
			uav_writeresponserequest => '0',                                                                                              --              (terminated)
			uav_writeresponsevalid   => open,                                                                                             --              (terminated)
			av_writeresponserequest  => open,                                                                                             --              (terminated)
			av_writeresponsevalid    => '0'                                                                                               --              (terminated)
		);

	capt3_0_avalon_parallel_port_slave_translator : component nios_system_ctr_moteur_avalon_parallel_port_slave_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 29,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 1,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 0,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => external_clocks_sys_clk_clk,                                                                   --                      clk.clk
			reset                    => cpu_jtag_debug_module_reset_reset,                                                             --                    reset.reset
			uav_address              => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => capt3_0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => capt3_0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => capt3_0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => capt3_0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => capt3_0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable            => capt3_0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_chipselect            => capt3_0_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_begintransfer         => open,                                                                                          --              (terminated)
			av_beginbursttransfer    => open,                                                                                          --              (terminated)
			av_burstcount            => open,                                                                                          --              (terminated)
			av_readdatavalid         => '0',                                                                                           --              (terminated)
			av_waitrequest           => '0',                                                                                           --              (terminated)
			av_writebyteenable       => open,                                                                                          --              (terminated)
			av_lock                  => open,                                                                                          --              (terminated)
			av_clken                 => open,                                                                                          --              (terminated)
			uav_clken                => '0',                                                                                           --              (terminated)
			av_debugaccess           => open,                                                                                          --              (terminated)
			av_outputenable          => open,                                                                                          --              (terminated)
			uav_response             => open,                                                                                          --              (terminated)
			av_response              => "00",                                                                                          --              (terminated)
			uav_writeresponserequest => '0',                                                                                           --              (terminated)
			uav_writeresponsevalid   => open,                                                                                          --              (terminated)
			av_writeresponserequest  => open,                                                                                          --              (terminated)
			av_writeresponsevalid    => '0'                                                                                            --              (terminated)
		);

	capt6_4_avalon_parallel_port_slave_translator : component nios_system_ctr_moteur_avalon_parallel_port_slave_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 29,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 1,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 0,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => external_clocks_sys_clk_clk,                                                                   --                      clk.clk
			reset                    => cpu_jtag_debug_module_reset_reset,                                                             --                    reset.reset
			uav_address              => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => capt6_4_avalon_parallel_port_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => capt6_4_avalon_parallel_port_slave_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => capt6_4_avalon_parallel_port_slave_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => capt6_4_avalon_parallel_port_slave_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => capt6_4_avalon_parallel_port_slave_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable            => capt6_4_avalon_parallel_port_slave_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_chipselect            => capt6_4_avalon_parallel_port_slave_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_begintransfer         => open,                                                                                          --              (terminated)
			av_beginbursttransfer    => open,                                                                                          --              (terminated)
			av_burstcount            => open,                                                                                          --              (terminated)
			av_readdatavalid         => '0',                                                                                           --              (terminated)
			av_waitrequest           => '0',                                                                                           --              (terminated)
			av_writebyteenable       => open,                                                                                          --              (terminated)
			av_lock                  => open,                                                                                          --              (terminated)
			av_clken                 => open,                                                                                          --              (terminated)
			uav_clken                => '0',                                                                                           --              (terminated)
			av_debugaccess           => open,                                                                                          --              (terminated)
			av_outputenable          => open,                                                                                          --              (terminated)
			uav_response             => open,                                                                                          --              (terminated)
			av_response              => "00",                                                                                          --              (terminated)
			uav_writeresponserequest => '0',                                                                                           --              (terminated)
			uav_writeresponsevalid   => open,                                                                                          --              (terminated)
			av_writeresponserequest  => open,                                                                                          --              (terminated)
			av_writeresponsevalid    => '0'                                                                                            --              (terminated)
		);

	cpu_instruction_master_translator_avalon_universal_master_0_agent : component altera_merlin_master_agent
		generic map (
			PKT_PROTECTION_H          => 95,
			PKT_PROTECTION_L          => 93,
			PKT_BEGIN_BURST           => 84,
			PKT_BURSTWRAP_H           => 76,
			PKT_BURSTWRAP_L           => 74,
			PKT_BURST_SIZE_H          => 79,
			PKT_BURST_SIZE_L          => 77,
			PKT_BURST_TYPE_H          => 81,
			PKT_BURST_TYPE_L          => 80,
			PKT_BYTE_CNT_H            => 73,
			PKT_BYTE_CNT_L            => 71,
			PKT_ADDR_H                => 64,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 65,
			PKT_TRANS_POSTED          => 66,
			PKT_TRANS_WRITE           => 67,
			PKT_TRANS_READ            => 68,
			PKT_TRANS_LOCK            => 69,
			PKT_TRANS_EXCLUSIVE       => 70,
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_SRC_ID_H              => 88,
			PKT_SRC_ID_L              => 86,
			PKT_DEST_ID_H             => 91,
			PKT_DEST_ID_L             => 89,
			PKT_THREAD_ID_H           => 92,
			PKT_THREAD_ID_L           => 92,
			PKT_CACHE_H               => 99,
			PKT_CACHE_L               => 96,
			PKT_DATA_SIDEBAND_H       => 83,
			PKT_DATA_SIDEBAND_L       => 83,
			PKT_QOS_H                 => 85,
			PKT_QOS_L                 => 85,
			PKT_ADDR_SIDEBAND_H       => 82,
			PKT_ADDR_SIDEBAND_L       => 82,
			PKT_RESPONSE_STATUS_H     => 101,
			PKT_RESPONSE_STATUS_L     => 100,
			ST_DATA_W                 => 102,
			ST_CHANNEL_W              => 8,
			AV_BURSTCOUNT_W           => 3,
			SUPPRESS_0_BYTEEN_RSP     => 0,
			ID                        => 1,
			BURSTWRAP_VALUE           => 3,
			CACHE_VALUE               => 0,
			SECURE_ACCESS_BIT         => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => external_clocks_sys_clk_clk,                                                        --       clk.clk
			reset                   => rst_controller_reset_out_reset,                                                     -- clk_reset.reset
			av_address              => cpu_instruction_master_translator_avalon_universal_master_0_address,                --        av.address
			av_write                => cpu_instruction_master_translator_avalon_universal_master_0_write,                  --          .write
			av_read                 => cpu_instruction_master_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata            => cpu_instruction_master_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata             => cpu_instruction_master_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest          => cpu_instruction_master_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid        => cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable           => cpu_instruction_master_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount           => cpu_instruction_master_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess          => cpu_instruction_master_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock                 => cpu_instruction_master_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid                => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data                 => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket        => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket          => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready                => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid                => limiter_rsp_src_valid,                                                              --        rp.valid
			rp_data                 => limiter_rsp_src_data,                                                               --          .data
			rp_channel              => limiter_rsp_src_channel,                                                            --          .channel
			rp_startofpacket        => limiter_rsp_src_startofpacket,                                                      --          .startofpacket
			rp_endofpacket          => limiter_rsp_src_endofpacket,                                                        --          .endofpacket
			rp_ready                => limiter_rsp_src_ready,                                                              --          .ready
			av_response             => open,                                                                               -- (terminated)
			av_writeresponserequest => '0',                                                                                -- (terminated)
			av_writeresponsevalid   => open                                                                                -- (terminated)
		);

	cpu_data_master_translator_avalon_universal_master_0_agent : component altera_merlin_master_agent
		generic map (
			PKT_PROTECTION_H          => 95,
			PKT_PROTECTION_L          => 93,
			PKT_BEGIN_BURST           => 84,
			PKT_BURSTWRAP_H           => 76,
			PKT_BURSTWRAP_L           => 74,
			PKT_BURST_SIZE_H          => 79,
			PKT_BURST_SIZE_L          => 77,
			PKT_BURST_TYPE_H          => 81,
			PKT_BURST_TYPE_L          => 80,
			PKT_BYTE_CNT_H            => 73,
			PKT_BYTE_CNT_L            => 71,
			PKT_ADDR_H                => 64,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 65,
			PKT_TRANS_POSTED          => 66,
			PKT_TRANS_WRITE           => 67,
			PKT_TRANS_READ            => 68,
			PKT_TRANS_LOCK            => 69,
			PKT_TRANS_EXCLUSIVE       => 70,
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_SRC_ID_H              => 88,
			PKT_SRC_ID_L              => 86,
			PKT_DEST_ID_H             => 91,
			PKT_DEST_ID_L             => 89,
			PKT_THREAD_ID_H           => 92,
			PKT_THREAD_ID_L           => 92,
			PKT_CACHE_H               => 99,
			PKT_CACHE_L               => 96,
			PKT_DATA_SIDEBAND_H       => 83,
			PKT_DATA_SIDEBAND_L       => 83,
			PKT_QOS_H                 => 85,
			PKT_QOS_L                 => 85,
			PKT_ADDR_SIDEBAND_H       => 82,
			PKT_ADDR_SIDEBAND_L       => 82,
			PKT_RESPONSE_STATUS_H     => 101,
			PKT_RESPONSE_STATUS_L     => 100,
			ST_DATA_W                 => 102,
			ST_CHANNEL_W              => 8,
			AV_BURSTCOUNT_W           => 3,
			SUPPRESS_0_BYTEEN_RSP     => 0,
			ID                        => 0,
			BURSTWRAP_VALUE           => 7,
			CACHE_VALUE               => 0,
			SECURE_ACCESS_BIT         => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => external_clocks_sys_clk_clk,                                                 --       clk.clk
			reset                   => rst_controller_reset_out_reset,                                              -- clk_reset.reset
			av_address              => cpu_data_master_translator_avalon_universal_master_0_address,                --        av.address
			av_write                => cpu_data_master_translator_avalon_universal_master_0_write,                  --          .write
			av_read                 => cpu_data_master_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata            => cpu_data_master_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata             => cpu_data_master_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest          => cpu_data_master_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid        => cpu_data_master_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable           => cpu_data_master_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount           => cpu_data_master_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess          => cpu_data_master_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock                 => cpu_data_master_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid                => cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data                 => cpu_data_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket        => cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket          => cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready                => cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid                => rsp_xbar_mux_001_src_valid,                                                  --        rp.valid
			rp_data                 => rsp_xbar_mux_001_src_data,                                                   --          .data
			rp_channel              => rsp_xbar_mux_001_src_channel,                                                --          .channel
			rp_startofpacket        => rsp_xbar_mux_001_src_startofpacket,                                          --          .startofpacket
			rp_endofpacket          => rsp_xbar_mux_001_src_endofpacket,                                            --          .endofpacket
			rp_ready                => rsp_xbar_mux_001_src_ready,                                                  --          .ready
			av_response             => open,                                                                        -- (terminated)
			av_writeresponserequest => '0',                                                                         -- (terminated)
			av_writeresponsevalid   => open                                                                         -- (terminated)
		);

	cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent : component nios_system_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 84,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 64,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 65,
			PKT_TRANS_POSTED          => 66,
			PKT_TRANS_WRITE           => 67,
			PKT_TRANS_READ            => 68,
			PKT_TRANS_LOCK            => 69,
			PKT_SRC_ID_H              => 88,
			PKT_SRC_ID_L              => 86,
			PKT_DEST_ID_H             => 91,
			PKT_DEST_ID_L             => 89,
			PKT_BURSTWRAP_H           => 76,
			PKT_BURSTWRAP_L           => 74,
			PKT_BYTE_CNT_H            => 73,
			PKT_BYTE_CNT_L            => 71,
			PKT_PROTECTION_H          => 95,
			PKT_PROTECTION_L          => 93,
			PKT_RESPONSE_STATUS_H     => 101,
			PKT_RESPONSE_STATUS_L     => 100,
			PKT_BURST_SIZE_H          => 79,
			PKT_BURST_SIZE_L          => 77,
			ST_CHANNEL_W              => 8,
			ST_DATA_W                 => 102,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => external_clocks_sys_clk_clk,                                                                --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                             --       clk_reset.reset
			m0_address              => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_src_ready,                                                                     --              cp.ready
			cp_valid                => cmd_xbar_mux_src_valid,                                                                     --                .valid
			cp_data                 => cmd_xbar_mux_src_data,                                                                      --                .data
			cp_startofpacket        => cmd_xbar_mux_src_startofpacket,                                                             --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_src_endofpacket,                                                               --                .endofpacket
			cp_channel              => cmd_xbar_mux_src_channel,                                                                   --                .channel
			rf_sink_ready           => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                       --     (terminated)
			m0_writeresponserequest => open,                                                                                       --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                         --     (terminated)
		);

	cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios_system_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 103,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => external_clocks_sys_clk_clk,                                                                --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                             -- clk_reset.reset
			in_data           => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                       -- (terminated)
			csr_read          => '0',                                                                                        -- (terminated)
			csr_write         => '0',                                                                                        -- (terminated)
			csr_readdata      => open,                                                                                       -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                         -- (terminated)
			almost_full_data  => open,                                                                                       -- (terminated)
			almost_empty_data => open,                                                                                       -- (terminated)
			in_empty          => '0',                                                                                        -- (terminated)
			out_empty         => open,                                                                                       -- (terminated)
			in_error          => '0',                                                                                        -- (terminated)
			out_error         => open,                                                                                       -- (terminated)
			in_channel        => '0',                                                                                        -- (terminated)
			out_channel       => open                                                                                        -- (terminated)
		);

	sdram_s1_translator_avalon_universal_slave_0_agent : component nios_system_sdram_s1_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 15,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 66,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 17,
			PKT_BYTEEN_L              => 16,
			PKT_ADDR_H                => 46,
			PKT_ADDR_L                => 18,
			PKT_TRANS_COMPRESSED_READ => 47,
			PKT_TRANS_POSTED          => 48,
			PKT_TRANS_WRITE           => 49,
			PKT_TRANS_READ            => 50,
			PKT_TRANS_LOCK            => 51,
			PKT_SRC_ID_H              => 70,
			PKT_SRC_ID_L              => 68,
			PKT_DEST_ID_H             => 73,
			PKT_DEST_ID_L             => 71,
			PKT_BURSTWRAP_H           => 58,
			PKT_BURSTWRAP_L           => 56,
			PKT_BYTE_CNT_H            => 55,
			PKT_BYTE_CNT_L            => 53,
			PKT_PROTECTION_H          => 77,
			PKT_PROTECTION_L          => 75,
			PKT_RESPONSE_STATUS_H     => 83,
			PKT_RESPONSE_STATUS_L     => 82,
			PKT_BURST_SIZE_H          => 61,
			PKT_BURST_SIZE_L          => 59,
			ST_CHANNEL_W              => 8,
			ST_DATA_W                 => 84,
			AVS_BURSTCOUNT_W          => 2,
			SUPPRESS_0_BYTEEN_CMD     => 1,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => external_clocks_sys_clk_clk,                                                   --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                --       clk_reset.reset
			m0_address              => sdram_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => sdram_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => sdram_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => sdram_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => burst_adapter_source0_ready,                                                   --              cp.ready
			cp_valid                => burst_adapter_source0_valid,                                                   --                .valid
			cp_data                 => burst_adapter_source0_data,                                                    --                .data
			cp_startofpacket        => burst_adapter_source0_startofpacket,                                           --                .startofpacket
			cp_endofpacket          => burst_adapter_source0_endofpacket,                                             --                .endofpacket
			cp_channel              => burst_adapter_source0_channel,                                                 --                .channel
			rf_sink_ready           => sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid,       --                .valid
			rdata_fifo_sink_data    => sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,        --                .data
			rdata_fifo_src_ready    => sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                          --     (terminated)
			m0_writeresponserequest => open,                                                                          --     (terminated)
			m0_writeresponsevalid   => '0'                                                                            --     (terminated)
		);

	sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios_system_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 85,
			FIFO_DEPTH          => 8,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => external_clocks_sys_clk_clk,                                                   --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                -- clk_reset.reset
			in_data           => sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                          -- (terminated)
			csr_read          => '0',                                                                           -- (terminated)
			csr_write         => '0',                                                                           -- (terminated)
			csr_readdata      => open,                                                                          -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                            -- (terminated)
			almost_full_data  => open,                                                                          -- (terminated)
			almost_empty_data => open,                                                                          -- (terminated)
			in_empty          => '0',                                                                           -- (terminated)
			out_empty         => open,                                                                          -- (terminated)
			in_error          => '0',                                                                           -- (terminated)
			out_error         => open,                                                                          -- (terminated)
			in_channel        => '0',                                                                           -- (terminated)
			out_channel       => open                                                                           -- (terminated)
		);

	sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo : component nios_system_sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 18,
			FIFO_DEPTH          => 8,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 0,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 3,
			USE_MEMORY_BLOCKS   => 1,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => external_clocks_sys_clk_clk,                                             --       clk.clk
			reset             => rst_controller_reset_out_reset,                                          -- clk_reset.reset
			in_data           => sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,  --        in.data
			in_valid          => sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid, --          .valid
			in_ready          => sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready, --          .ready
			out_data          => sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,  --       out.data
			out_valid         => sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid, --          .valid
			out_ready         => sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready, --          .ready
			csr_address       => "00",                                                                    -- (terminated)
			csr_read          => '0',                                                                     -- (terminated)
			csr_write         => '0',                                                                     -- (terminated)
			csr_readdata      => open,                                                                    -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                      -- (terminated)
			almost_full_data  => open,                                                                    -- (terminated)
			almost_empty_data => open,                                                                    -- (terminated)
			in_startofpacket  => '0',                                                                     -- (terminated)
			in_endofpacket    => '0',                                                                     -- (terminated)
			out_startofpacket => open,                                                                    -- (terminated)
			out_endofpacket   => open,                                                                    -- (terminated)
			in_empty          => '0',                                                                     -- (terminated)
			out_empty         => open,                                                                    -- (terminated)
			in_error          => '0',                                                                     -- (terminated)
			out_error         => open,                                                                    -- (terminated)
			in_channel        => '0',                                                                     -- (terminated)
			out_channel       => open                                                                     -- (terminated)
		);

	interval_timer_s1_translator_avalon_universal_slave_0_agent : component nios_system_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 84,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 64,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 65,
			PKT_TRANS_POSTED          => 66,
			PKT_TRANS_WRITE           => 67,
			PKT_TRANS_READ            => 68,
			PKT_TRANS_LOCK            => 69,
			PKT_SRC_ID_H              => 88,
			PKT_SRC_ID_L              => 86,
			PKT_DEST_ID_H             => 91,
			PKT_DEST_ID_L             => 89,
			PKT_BURSTWRAP_H           => 76,
			PKT_BURSTWRAP_L           => 74,
			PKT_BYTE_CNT_H            => 73,
			PKT_BYTE_CNT_L            => 71,
			PKT_PROTECTION_H          => 95,
			PKT_PROTECTION_L          => 93,
			PKT_RESPONSE_STATUS_H     => 101,
			PKT_RESPONSE_STATUS_L     => 100,
			PKT_BURST_SIZE_H          => 79,
			PKT_BURST_SIZE_L          => 77,
			ST_CHANNEL_W              => 8,
			ST_DATA_W                 => 102,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => external_clocks_sys_clk_clk,                                                            --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                         --       clk_reset.reset
			m0_address              => interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => interval_timer_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src2_ready,                                                          --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src2_valid,                                                          --                .valid
			cp_data                 => cmd_xbar_demux_001_src2_data,                                                           --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src2_startofpacket,                                                  --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src2_endofpacket,                                                    --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src2_channel,                                                        --                .channel
			rf_sink_ready           => interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => interval_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => interval_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => interval_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => interval_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => interval_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => interval_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                   --     (terminated)
			m0_writeresponserequest => open,                                                                                   --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                     --     (terminated)
		);

	interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios_system_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 103,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => external_clocks_sys_clk_clk,                                                            --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                         -- clk_reset.reset
			in_data           => interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => interval_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => interval_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                   -- (terminated)
			csr_read          => '0',                                                                                    -- (terminated)
			csr_write         => '0',                                                                                    -- (terminated)
			csr_readdata      => open,                                                                                   -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                     -- (terminated)
			almost_full_data  => open,                                                                                   -- (terminated)
			almost_empty_data => open,                                                                                   -- (terminated)
			in_empty          => '0',                                                                                    -- (terminated)
			out_empty         => open,                                                                                   -- (terminated)
			in_error          => '0',                                                                                    -- (terminated)
			out_error         => open,                                                                                   -- (terminated)
			in_channel        => '0',                                                                                    -- (terminated)
			out_channel       => open                                                                                    -- (terminated)
		);

	sysid_control_slave_translator_avalon_universal_slave_0_agent : component nios_system_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 84,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 64,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 65,
			PKT_TRANS_POSTED          => 66,
			PKT_TRANS_WRITE           => 67,
			PKT_TRANS_READ            => 68,
			PKT_TRANS_LOCK            => 69,
			PKT_SRC_ID_H              => 88,
			PKT_SRC_ID_L              => 86,
			PKT_DEST_ID_H             => 91,
			PKT_DEST_ID_L             => 89,
			PKT_BURSTWRAP_H           => 76,
			PKT_BURSTWRAP_L           => 74,
			PKT_BYTE_CNT_H            => 73,
			PKT_BYTE_CNT_L            => 71,
			PKT_PROTECTION_H          => 95,
			PKT_PROTECTION_L          => 93,
			PKT_RESPONSE_STATUS_H     => 101,
			PKT_RESPONSE_STATUS_L     => 100,
			PKT_BURST_SIZE_H          => 79,
			PKT_BURST_SIZE_L          => 77,
			ST_CHANNEL_W              => 8,
			ST_DATA_W                 => 102,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => external_clocks_sys_clk_clk,                                                              --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                           --       clk_reset.reset
			m0_address              => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src3_ready,                                                            --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src3_valid,                                                            --                .valid
			cp_data                 => cmd_xbar_demux_001_src3_data,                                                             --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src3_startofpacket,                                                    --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src3_endofpacket,                                                      --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src3_channel,                                                          --                .channel
			rf_sink_ready           => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                     --     (terminated)
			m0_writeresponserequest => open,                                                                                     --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                       --     (terminated)
		);

	sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios_system_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 103,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => external_clocks_sys_clk_clk,                                                              --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                           -- clk_reset.reset
			in_data           => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                     -- (terminated)
			csr_read          => '0',                                                                                      -- (terminated)
			csr_write         => '0',                                                                                      -- (terminated)
			csr_readdata      => open,                                                                                     -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                       -- (terminated)
			almost_full_data  => open,                                                                                     -- (terminated)
			almost_empty_data => open,                                                                                     -- (terminated)
			in_empty          => '0',                                                                                      -- (terminated)
			out_empty         => open,                                                                                     -- (terminated)
			in_error          => '0',                                                                                      -- (terminated)
			out_error         => open,                                                                                     -- (terminated)
			in_channel        => '0',                                                                                      -- (terminated)
			out_channel       => open                                                                                      -- (terminated)
		);

	jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent : component nios_system_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 84,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 64,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 65,
			PKT_TRANS_POSTED          => 66,
			PKT_TRANS_WRITE           => 67,
			PKT_TRANS_READ            => 68,
			PKT_TRANS_LOCK            => 69,
			PKT_SRC_ID_H              => 88,
			PKT_SRC_ID_L              => 86,
			PKT_DEST_ID_H             => 91,
			PKT_DEST_ID_L             => 89,
			PKT_BURSTWRAP_H           => 76,
			PKT_BURSTWRAP_L           => 74,
			PKT_BYTE_CNT_H            => 73,
			PKT_BYTE_CNT_L            => 71,
			PKT_PROTECTION_H          => 95,
			PKT_PROTECTION_L          => 93,
			PKT_RESPONSE_STATUS_H     => 101,
			PKT_RESPONSE_STATUS_L     => 100,
			PKT_BURST_SIZE_H          => 79,
			PKT_BURST_SIZE_L          => 77,
			ST_CHANNEL_W              => 8,
			ST_DATA_W                 => 102,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => external_clocks_sys_clk_clk,                                                                      --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                                   --       clk_reset.reset
			m0_address              => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src4_ready,                                                                    --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src4_valid,                                                                    --                .valid
			cp_data                 => cmd_xbar_demux_001_src4_data,                                                                     --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src4_startofpacket,                                                            --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src4_endofpacket,                                                              --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src4_channel,                                                                  --                .channel
			rf_sink_ready           => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                             --     (terminated)
			m0_writeresponserequest => open,                                                                                             --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                               --     (terminated)
		);

	jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios_system_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 103,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => external_clocks_sys_clk_clk,                                                                      --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                                   -- clk_reset.reset
			in_data           => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                             -- (terminated)
			csr_read          => '0',                                                                                              -- (terminated)
			csr_write         => '0',                                                                                              -- (terminated)
			csr_readdata      => open,                                                                                             -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                               -- (terminated)
			almost_full_data  => open,                                                                                             -- (terminated)
			almost_empty_data => open,                                                                                             -- (terminated)
			in_empty          => '0',                                                                                              -- (terminated)
			out_empty         => open,                                                                                             -- (terminated)
			in_error          => '0',                                                                                              -- (terminated)
			out_error         => open,                                                                                             -- (terminated)
			in_channel        => '0',                                                                                              -- (terminated)
			out_channel       => open                                                                                              -- (terminated)
		);

	ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent : component nios_system_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 84,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 64,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 65,
			PKT_TRANS_POSTED          => 66,
			PKT_TRANS_WRITE           => 67,
			PKT_TRANS_READ            => 68,
			PKT_TRANS_LOCK            => 69,
			PKT_SRC_ID_H              => 88,
			PKT_SRC_ID_L              => 86,
			PKT_DEST_ID_H             => 91,
			PKT_DEST_ID_L             => 89,
			PKT_BURSTWRAP_H           => 76,
			PKT_BURSTWRAP_L           => 74,
			PKT_BYTE_CNT_H            => 73,
			PKT_BYTE_CNT_L            => 71,
			PKT_PROTECTION_H          => 95,
			PKT_PROTECTION_L          => 93,
			PKT_RESPONSE_STATUS_H     => 101,
			PKT_RESPONSE_STATUS_L     => 100,
			PKT_BURST_SIZE_H          => 79,
			PKT_BURST_SIZE_L          => 77,
			ST_CHANNEL_W              => 8,
			ST_DATA_W                 => 102,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => external_clocks_sys_clk_clk,                                                                                --             clk.clk
			reset                   => cpu_jtag_debug_module_reset_reset,                                                                          --       clk_reset.reset
			m0_address              => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src5_ready,                                                                              --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src5_valid,                                                                              --                .valid
			cp_data                 => cmd_xbar_demux_001_src5_data,                                                                               --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src5_startofpacket,                                                                      --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src5_endofpacket,                                                                        --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src5_channel,                                                                            --                .channel
			rf_sink_ready           => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                                       --     (terminated)
			m0_writeresponserequest => open,                                                                                                       --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                                         --     (terminated)
		);

	ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios_system_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 103,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => external_clocks_sys_clk_clk,                                                                                --       clk.clk
			reset             => cpu_jtag_debug_module_reset_reset,                                                                          -- clk_reset.reset
			in_data           => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                                       -- (terminated)
			csr_read          => '0',                                                                                                        -- (terminated)
			csr_write         => '0',                                                                                                        -- (terminated)
			csr_readdata      => open,                                                                                                       -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                                         -- (terminated)
			almost_full_data  => open,                                                                                                       -- (terminated)
			almost_empty_data => open,                                                                                                       -- (terminated)
			in_empty          => '0',                                                                                                        -- (terminated)
			out_empty         => open,                                                                                                       -- (terminated)
			in_error          => '0',                                                                                                        -- (terminated)
			out_error         => open,                                                                                                       -- (terminated)
			in_channel        => '0',                                                                                                        -- (terminated)
			out_channel       => open                                                                                                        -- (terminated)
		);

	capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent : component nios_system_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 84,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 64,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 65,
			PKT_TRANS_POSTED          => 66,
			PKT_TRANS_WRITE           => 67,
			PKT_TRANS_READ            => 68,
			PKT_TRANS_LOCK            => 69,
			PKT_SRC_ID_H              => 88,
			PKT_SRC_ID_L              => 86,
			PKT_DEST_ID_H             => 91,
			PKT_DEST_ID_L             => 89,
			PKT_BURSTWRAP_H           => 76,
			PKT_BURSTWRAP_L           => 74,
			PKT_BYTE_CNT_H            => 73,
			PKT_BYTE_CNT_L            => 71,
			PKT_PROTECTION_H          => 95,
			PKT_PROTECTION_L          => 93,
			PKT_RESPONSE_STATUS_H     => 101,
			PKT_RESPONSE_STATUS_L     => 100,
			PKT_BURST_SIZE_H          => 79,
			PKT_BURST_SIZE_L          => 77,
			ST_CHANNEL_W              => 8,
			ST_DATA_W                 => 102,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => external_clocks_sys_clk_clk,                                                                             --             clk.clk
			reset                   => cpu_jtag_debug_module_reset_reset,                                                                       --       clk_reset.reset
			m0_address              => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src6_ready,                                                                           --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src6_valid,                                                                           --                .valid
			cp_data                 => cmd_xbar_demux_001_src6_data,                                                                            --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src6_startofpacket,                                                                   --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src6_endofpacket,                                                                     --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src6_channel,                                                                         --                .channel
			rf_sink_ready           => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                                    --     (terminated)
			m0_writeresponserequest => open,                                                                                                    --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                                      --     (terminated)
		);

	capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios_system_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 103,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => external_clocks_sys_clk_clk,                                                                             --       clk.clk
			reset             => cpu_jtag_debug_module_reset_reset,                                                                       -- clk_reset.reset
			in_data           => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                                    -- (terminated)
			csr_read          => '0',                                                                                                     -- (terminated)
			csr_write         => '0',                                                                                                     -- (terminated)
			csr_readdata      => open,                                                                                                    -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                                      -- (terminated)
			almost_full_data  => open,                                                                                                    -- (terminated)
			almost_empty_data => open,                                                                                                    -- (terminated)
			in_empty          => '0',                                                                                                     -- (terminated)
			out_empty         => open,                                                                                                    -- (terminated)
			in_error          => '0',                                                                                                     -- (terminated)
			out_error         => open,                                                                                                    -- (terminated)
			in_channel        => '0',                                                                                                     -- (terminated)
			out_channel       => open                                                                                                     -- (terminated)
		);

	capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent : component nios_system_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 84,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 64,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 65,
			PKT_TRANS_POSTED          => 66,
			PKT_TRANS_WRITE           => 67,
			PKT_TRANS_READ            => 68,
			PKT_TRANS_LOCK            => 69,
			PKT_SRC_ID_H              => 88,
			PKT_SRC_ID_L              => 86,
			PKT_DEST_ID_H             => 91,
			PKT_DEST_ID_L             => 89,
			PKT_BURSTWRAP_H           => 76,
			PKT_BURSTWRAP_L           => 74,
			PKT_BYTE_CNT_H            => 73,
			PKT_BYTE_CNT_L            => 71,
			PKT_PROTECTION_H          => 95,
			PKT_PROTECTION_L          => 93,
			PKT_RESPONSE_STATUS_H     => 101,
			PKT_RESPONSE_STATUS_L     => 100,
			PKT_BURST_SIZE_H          => 79,
			PKT_BURST_SIZE_L          => 77,
			ST_CHANNEL_W              => 8,
			ST_DATA_W                 => 102,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => external_clocks_sys_clk_clk,                                                                             --             clk.clk
			reset                   => cpu_jtag_debug_module_reset_reset,                                                                       --       clk_reset.reset
			m0_address              => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src7_ready,                                                                           --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src7_valid,                                                                           --                .valid
			cp_data                 => cmd_xbar_demux_001_src7_data,                                                                            --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src7_startofpacket,                                                                   --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src7_endofpacket,                                                                     --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src7_channel,                                                                         --                .channel
			rf_sink_ready           => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                                    --     (terminated)
			m0_writeresponserequest => open,                                                                                                    --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                                      --     (terminated)
		);

	capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios_system_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 103,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => external_clocks_sys_clk_clk,                                                                             --       clk.clk
			reset             => cpu_jtag_debug_module_reset_reset,                                                                       -- clk_reset.reset
			in_data           => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                                    -- (terminated)
			csr_read          => '0',                                                                                                     -- (terminated)
			csr_write         => '0',                                                                                                     -- (terminated)
			csr_readdata      => open,                                                                                                    -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                                      -- (terminated)
			almost_full_data  => open,                                                                                                    -- (terminated)
			almost_empty_data => open,                                                                                                    -- (terminated)
			in_empty          => '0',                                                                                                     -- (terminated)
			out_empty         => open,                                                                                                    -- (terminated)
			in_error          => '0',                                                                                                     -- (terminated)
			out_error         => open,                                                                                                    -- (terminated)
			in_channel        => '0',                                                                                                     -- (terminated)
			out_channel       => open                                                                                                     -- (terminated)
		);

	addr_router : component nios_system_addr_router
		port map (
			sink_ready         => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => external_clocks_sys_clk_clk,                                                        --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                     -- clk_reset.reset
			src_ready          => addr_router_src_ready,                                                              --       src.ready
			src_valid          => addr_router_src_valid,                                                              --          .valid
			src_data           => addr_router_src_data,                                                               --          .data
			src_channel        => addr_router_src_channel,                                                            --          .channel
			src_startofpacket  => addr_router_src_startofpacket,                                                      --          .startofpacket
			src_endofpacket    => addr_router_src_endofpacket                                                         --          .endofpacket
		);

	addr_router_001 : component nios_system_addr_router_001
		port map (
			sink_ready         => cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => cpu_data_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => external_clocks_sys_clk_clk,                                                 --       clk.clk
			reset              => rst_controller_reset_out_reset,                                              -- clk_reset.reset
			src_ready          => addr_router_001_src_ready,                                                   --       src.ready
			src_valid          => addr_router_001_src_valid,                                                   --          .valid
			src_data           => addr_router_001_src_data,                                                    --          .data
			src_channel        => addr_router_001_src_channel,                                                 --          .channel
			src_startofpacket  => addr_router_001_src_startofpacket,                                           --          .startofpacket
			src_endofpacket    => addr_router_001_src_endofpacket                                              --          .endofpacket
		);

	id_router : component nios_system_id_router
		port map (
			sink_ready         => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => external_clocks_sys_clk_clk,                                                      --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                   -- clk_reset.reset
			src_ready          => id_router_src_ready,                                                              --       src.ready
			src_valid          => id_router_src_valid,                                                              --          .valid
			src_data           => id_router_src_data,                                                               --          .data
			src_channel        => id_router_src_channel,                                                            --          .channel
			src_startofpacket  => id_router_src_startofpacket,                                                      --          .startofpacket
			src_endofpacket    => id_router_src_endofpacket                                                         --          .endofpacket
		);

	id_router_001 : component nios_system_id_router_001
		port map (
			sink_ready         => sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => sdram_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => external_clocks_sys_clk_clk,                                         --       clk.clk
			reset              => rst_controller_reset_out_reset,                                      -- clk_reset.reset
			src_ready          => id_router_001_src_ready,                                             --       src.ready
			src_valid          => id_router_001_src_valid,                                             --          .valid
			src_data           => id_router_001_src_data,                                              --          .data
			src_channel        => id_router_001_src_channel,                                           --          .channel
			src_startofpacket  => id_router_001_src_startofpacket,                                     --          .startofpacket
			src_endofpacket    => id_router_001_src_endofpacket                                        --          .endofpacket
		);

	id_router_002 : component nios_system_id_router_002
		port map (
			sink_ready         => interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => interval_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => external_clocks_sys_clk_clk,                                                  --       clk.clk
			reset              => rst_controller_reset_out_reset,                                               -- clk_reset.reset
			src_ready          => id_router_002_src_ready,                                                      --       src.ready
			src_valid          => id_router_002_src_valid,                                                      --          .valid
			src_data           => id_router_002_src_data,                                                       --          .data
			src_channel        => id_router_002_src_channel,                                                    --          .channel
			src_startofpacket  => id_router_002_src_startofpacket,                                              --          .startofpacket
			src_endofpacket    => id_router_002_src_endofpacket                                                 --          .endofpacket
		);

	id_router_003 : component nios_system_id_router_002
		port map (
			sink_ready         => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => external_clocks_sys_clk_clk,                                                    --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                 -- clk_reset.reset
			src_ready          => id_router_003_src_ready,                                                        --       src.ready
			src_valid          => id_router_003_src_valid,                                                        --          .valid
			src_data           => id_router_003_src_data,                                                         --          .data
			src_channel        => id_router_003_src_channel,                                                      --          .channel
			src_startofpacket  => id_router_003_src_startofpacket,                                                --          .startofpacket
			src_endofpacket    => id_router_003_src_endofpacket                                                   --          .endofpacket
		);

	id_router_004 : component nios_system_id_router_002
		port map (
			sink_ready         => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => external_clocks_sys_clk_clk,                                                            --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                         -- clk_reset.reset
			src_ready          => id_router_004_src_ready,                                                                --       src.ready
			src_valid          => id_router_004_src_valid,                                                                --          .valid
			src_data           => id_router_004_src_data,                                                                 --          .data
			src_channel        => id_router_004_src_channel,                                                              --          .channel
			src_startofpacket  => id_router_004_src_startofpacket,                                                        --          .startofpacket
			src_endofpacket    => id_router_004_src_endofpacket                                                           --          .endofpacket
		);

	id_router_005 : component nios_system_id_router_002
		port map (
			sink_ready         => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => ctr_moteur_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => external_clocks_sys_clk_clk,                                                                      --       clk.clk
			reset              => cpu_jtag_debug_module_reset_reset,                                                                -- clk_reset.reset
			src_ready          => id_router_005_src_ready,                                                                          --       src.ready
			src_valid          => id_router_005_src_valid,                                                                          --          .valid
			src_data           => id_router_005_src_data,                                                                           --          .data
			src_channel        => id_router_005_src_channel,                                                                        --          .channel
			src_startofpacket  => id_router_005_src_startofpacket,                                                                  --          .startofpacket
			src_endofpacket    => id_router_005_src_endofpacket                                                                     --          .endofpacket
		);

	id_router_006 : component nios_system_id_router_002
		port map (
			sink_ready         => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => capt3_0_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => external_clocks_sys_clk_clk,                                                                   --       clk.clk
			reset              => cpu_jtag_debug_module_reset_reset,                                                             -- clk_reset.reset
			src_ready          => id_router_006_src_ready,                                                                       --       src.ready
			src_valid          => id_router_006_src_valid,                                                                       --          .valid
			src_data           => id_router_006_src_data,                                                                        --          .data
			src_channel        => id_router_006_src_channel,                                                                     --          .channel
			src_startofpacket  => id_router_006_src_startofpacket,                                                               --          .startofpacket
			src_endofpacket    => id_router_006_src_endofpacket                                                                  --          .endofpacket
		);

	id_router_007 : component nios_system_id_router_002
		port map (
			sink_ready         => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => capt6_4_avalon_parallel_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => external_clocks_sys_clk_clk,                                                                   --       clk.clk
			reset              => cpu_jtag_debug_module_reset_reset,                                                             -- clk_reset.reset
			src_ready          => id_router_007_src_ready,                                                                       --       src.ready
			src_valid          => id_router_007_src_valid,                                                                       --          .valid
			src_data           => id_router_007_src_data,                                                                        --          .data
			src_channel        => id_router_007_src_channel,                                                                     --          .channel
			src_startofpacket  => id_router_007_src_startofpacket,                                                               --          .startofpacket
			src_endofpacket    => id_router_007_src_endofpacket                                                                  --          .endofpacket
		);

	limiter : component altera_merlin_traffic_limiter
		generic map (
			PKT_DEST_ID_H             => 91,
			PKT_DEST_ID_L             => 89,
			PKT_TRANS_POSTED          => 66,
			PKT_TRANS_WRITE           => 67,
			MAX_OUTSTANDING_RESPONSES => 9,
			PIPELINED                 => 0,
			ST_DATA_W                 => 102,
			ST_CHANNEL_W              => 8,
			VALID_WIDTH               => 8,
			ENFORCE_ORDER             => 1,
			PREVENT_HAZARDS           => 0,
			PKT_BYTE_CNT_H            => 73,
			PKT_BYTE_CNT_L            => 71,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32
		)
		port map (
			clk                    => external_clocks_sys_clk_clk,    --       clk.clk
			reset                  => rst_controller_reset_out_reset, -- clk_reset.reset
			cmd_sink_ready         => addr_router_src_ready,          --  cmd_sink.ready
			cmd_sink_valid         => addr_router_src_valid,          --          .valid
			cmd_sink_data          => addr_router_src_data,           --          .data
			cmd_sink_channel       => addr_router_src_channel,        --          .channel
			cmd_sink_startofpacket => addr_router_src_startofpacket,  --          .startofpacket
			cmd_sink_endofpacket   => addr_router_src_endofpacket,    --          .endofpacket
			cmd_src_ready          => limiter_cmd_src_ready,          --   cmd_src.ready
			cmd_src_data           => limiter_cmd_src_data,           --          .data
			cmd_src_channel        => limiter_cmd_src_channel,        --          .channel
			cmd_src_startofpacket  => limiter_cmd_src_startofpacket,  --          .startofpacket
			cmd_src_endofpacket    => limiter_cmd_src_endofpacket,    --          .endofpacket
			rsp_sink_ready         => rsp_xbar_mux_src_ready,         --  rsp_sink.ready
			rsp_sink_valid         => rsp_xbar_mux_src_valid,         --          .valid
			rsp_sink_channel       => rsp_xbar_mux_src_channel,       --          .channel
			rsp_sink_data          => rsp_xbar_mux_src_data,          --          .data
			rsp_sink_startofpacket => rsp_xbar_mux_src_startofpacket, --          .startofpacket
			rsp_sink_endofpacket   => rsp_xbar_mux_src_endofpacket,   --          .endofpacket
			rsp_src_ready          => limiter_rsp_src_ready,          --   rsp_src.ready
			rsp_src_valid          => limiter_rsp_src_valid,          --          .valid
			rsp_src_data           => limiter_rsp_src_data,           --          .data
			rsp_src_channel        => limiter_rsp_src_channel,        --          .channel
			rsp_src_startofpacket  => limiter_rsp_src_startofpacket,  --          .startofpacket
			rsp_src_endofpacket    => limiter_rsp_src_endofpacket,    --          .endofpacket
			cmd_src_valid          => limiter_cmd_valid_data          -- cmd_valid.data
		);

	burst_adapter : component altera_merlin_burst_adapter
		generic map (
			PKT_ADDR_H                => 46,
			PKT_ADDR_L                => 18,
			PKT_BEGIN_BURST           => 66,
			PKT_BYTE_CNT_H            => 55,
			PKT_BYTE_CNT_L            => 53,
			PKT_BYTEEN_H              => 17,
			PKT_BYTEEN_L              => 16,
			PKT_BURST_SIZE_H          => 61,
			PKT_BURST_SIZE_L          => 59,
			PKT_BURST_TYPE_H          => 63,
			PKT_BURST_TYPE_L          => 62,
			PKT_BURSTWRAP_H           => 58,
			PKT_BURSTWRAP_L           => 56,
			PKT_TRANS_COMPRESSED_READ => 47,
			PKT_TRANS_WRITE           => 49,
			PKT_TRANS_READ            => 50,
			OUT_NARROW_SIZE           => 0,
			IN_NARROW_SIZE            => 0,
			OUT_FIXED                 => 0,
			OUT_COMPLETE_WRAP         => 0,
			ST_DATA_W                 => 84,
			ST_CHANNEL_W              => 8,
			OUT_BYTE_CNT_H            => 54,
			OUT_BURSTWRAP_H           => 58,
			COMPRESSED_READ_SUPPORT   => 0,
			BYTEENABLE_SYNTHESIS      => 1,
			PIPE_INPUTS               => 0,
			NO_WRAP_SUPPORT           => 0,
			BURSTWRAP_CONST_MASK      => 3,
			BURSTWRAP_CONST_VALUE     => 3
		)
		port map (
			clk                   => external_clocks_sys_clk_clk,         --       cr0.clk
			reset                 => rst_controller_reset_out_reset,      -- cr0_reset.reset
			sink0_valid           => width_adapter_src_valid,             --     sink0.valid
			sink0_data            => width_adapter_src_data,              --          .data
			sink0_channel         => width_adapter_src_channel,           --          .channel
			sink0_startofpacket   => width_adapter_src_startofpacket,     --          .startofpacket
			sink0_endofpacket     => width_adapter_src_endofpacket,       --          .endofpacket
			sink0_ready           => width_adapter_src_ready,             --          .ready
			source0_valid         => burst_adapter_source0_valid,         --   source0.valid
			source0_data          => burst_adapter_source0_data,          --          .data
			source0_channel       => burst_adapter_source0_channel,       --          .channel
			source0_startofpacket => burst_adapter_source0_startofpacket, --          .startofpacket
			source0_endofpacket   => burst_adapter_source0_endofpacket,   --          .endofpacket
			source0_ready         => burst_adapter_source0_ready          --          .ready
		);

	rst_controller : component nios_system_rst_controller
		generic map (
			NUM_RESET_INPUTS        => 2,
			OUTPUT_RESET_SYNC_EDGES => "deassert",
			SYNC_DEPTH              => 2,
			RESET_REQUEST_PRESENT   => 0
		)
		port map (
			reset_in0  => reset_n_ports_inv,                 -- reset_in0.reset
			reset_in1  => cpu_jtag_debug_module_reset_reset, -- reset_in1.reset
			clk        => external_clocks_sys_clk_clk,       --       clk.clk
			reset_out  => rst_controller_reset_out_reset,    -- reset_out.reset
			reset_req  => open,                              -- (terminated)
			reset_in2  => '0',                               -- (terminated)
			reset_in3  => '0',                               -- (terminated)
			reset_in4  => '0',                               -- (terminated)
			reset_in5  => '0',                               -- (terminated)
			reset_in6  => '0',                               -- (terminated)
			reset_in7  => '0',                               -- (terminated)
			reset_in8  => '0',                               -- (terminated)
			reset_in9  => '0',                               -- (terminated)
			reset_in10 => '0',                               -- (terminated)
			reset_in11 => '0',                               -- (terminated)
			reset_in12 => '0',                               -- (terminated)
			reset_in13 => '0',                               -- (terminated)
			reset_in14 => '0',                               -- (terminated)
			reset_in15 => '0'                                -- (terminated)
		);

	rst_controller_001 : component nios_system_rst_controller_001
		generic map (
			NUM_RESET_INPUTS        => 1,
			OUTPUT_RESET_SYNC_EDGES => "deassert",
			SYNC_DEPTH              => 2,
			RESET_REQUEST_PRESENT   => 0
		)
		port map (
			reset_in0  => reset_n_ports_inv,                  -- reset_in0.reset
			clk        => clk,                                --       clk.clk
			reset_out  => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req  => open,                               -- (terminated)
			reset_in1  => '0',                                -- (terminated)
			reset_in2  => '0',                                -- (terminated)
			reset_in3  => '0',                                -- (terminated)
			reset_in4  => '0',                                -- (terminated)
			reset_in5  => '0',                                -- (terminated)
			reset_in6  => '0',                                -- (terminated)
			reset_in7  => '0',                                -- (terminated)
			reset_in8  => '0',                                -- (terminated)
			reset_in9  => '0',                                -- (terminated)
			reset_in10 => '0',                                -- (terminated)
			reset_in11 => '0',                                -- (terminated)
			reset_in12 => '0',                                -- (terminated)
			reset_in13 => '0',                                -- (terminated)
			reset_in14 => '0',                                -- (terminated)
			reset_in15 => '0'                                 -- (terminated)
		);

	cmd_xbar_demux : component nios_system_cmd_xbar_demux
		port map (
			clk                => external_clocks_sys_clk_clk,       --        clk.clk
			reset              => rst_controller_reset_out_reset,    --  clk_reset.reset
			sink_ready         => limiter_cmd_src_ready,             --       sink.ready
			sink_channel       => limiter_cmd_src_channel,           --           .channel
			sink_data          => limiter_cmd_src_data,              --           .data
			sink_startofpacket => limiter_cmd_src_startofpacket,     --           .startofpacket
			sink_endofpacket   => limiter_cmd_src_endofpacket,       --           .endofpacket
			sink_valid         => limiter_cmd_valid_data,            -- sink_valid.data
			src0_ready         => cmd_xbar_demux_src0_ready,         --       src0.ready
			src0_valid         => cmd_xbar_demux_src0_valid,         --           .valid
			src0_data          => cmd_xbar_demux_src0_data,          --           .data
			src0_channel       => cmd_xbar_demux_src0_channel,       --           .channel
			src0_startofpacket => cmd_xbar_demux_src0_startofpacket, --           .startofpacket
			src0_endofpacket   => cmd_xbar_demux_src0_endofpacket,   --           .endofpacket
			src1_ready         => cmd_xbar_demux_src1_ready,         --       src1.ready
			src1_valid         => cmd_xbar_demux_src1_valid,         --           .valid
			src1_data          => cmd_xbar_demux_src1_data,          --           .data
			src1_channel       => cmd_xbar_demux_src1_channel,       --           .channel
			src1_startofpacket => cmd_xbar_demux_src1_startofpacket, --           .startofpacket
			src1_endofpacket   => cmd_xbar_demux_src1_endofpacket    --           .endofpacket
		);

	cmd_xbar_demux_001 : component nios_system_cmd_xbar_demux_001
		port map (
			clk                => external_clocks_sys_clk_clk,           --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => addr_router_001_src_ready,             --      sink.ready
			sink_channel       => addr_router_001_src_channel,           --          .channel
			sink_data          => addr_router_001_src_data,              --          .data
			sink_startofpacket => addr_router_001_src_startofpacket,     --          .startofpacket
			sink_endofpacket   => addr_router_001_src_endofpacket,       --          .endofpacket
			sink_valid(0)      => addr_router_001_src_valid,             --          .valid
			src0_ready         => cmd_xbar_demux_001_src0_ready,         --      src0.ready
			src0_valid         => cmd_xbar_demux_001_src0_valid,         --          .valid
			src0_data          => cmd_xbar_demux_001_src0_data,          --          .data
			src0_channel       => cmd_xbar_demux_001_src0_channel,       --          .channel
			src0_startofpacket => cmd_xbar_demux_001_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => cmd_xbar_demux_001_src0_endofpacket,   --          .endofpacket
			src1_ready         => cmd_xbar_demux_001_src1_ready,         --      src1.ready
			src1_valid         => cmd_xbar_demux_001_src1_valid,         --          .valid
			src1_data          => cmd_xbar_demux_001_src1_data,          --          .data
			src1_channel       => cmd_xbar_demux_001_src1_channel,       --          .channel
			src1_startofpacket => cmd_xbar_demux_001_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => cmd_xbar_demux_001_src1_endofpacket,   --          .endofpacket
			src2_ready         => cmd_xbar_demux_001_src2_ready,         --      src2.ready
			src2_valid         => cmd_xbar_demux_001_src2_valid,         --          .valid
			src2_data          => cmd_xbar_demux_001_src2_data,          --          .data
			src2_channel       => cmd_xbar_demux_001_src2_channel,       --          .channel
			src2_startofpacket => cmd_xbar_demux_001_src2_startofpacket, --          .startofpacket
			src2_endofpacket   => cmd_xbar_demux_001_src2_endofpacket,   --          .endofpacket
			src3_ready         => cmd_xbar_demux_001_src3_ready,         --      src3.ready
			src3_valid         => cmd_xbar_demux_001_src3_valid,         --          .valid
			src3_data          => cmd_xbar_demux_001_src3_data,          --          .data
			src3_channel       => cmd_xbar_demux_001_src3_channel,       --          .channel
			src3_startofpacket => cmd_xbar_demux_001_src3_startofpacket, --          .startofpacket
			src3_endofpacket   => cmd_xbar_demux_001_src3_endofpacket,   --          .endofpacket
			src4_ready         => cmd_xbar_demux_001_src4_ready,         --      src4.ready
			src4_valid         => cmd_xbar_demux_001_src4_valid,         --          .valid
			src4_data          => cmd_xbar_demux_001_src4_data,          --          .data
			src4_channel       => cmd_xbar_demux_001_src4_channel,       --          .channel
			src4_startofpacket => cmd_xbar_demux_001_src4_startofpacket, --          .startofpacket
			src4_endofpacket   => cmd_xbar_demux_001_src4_endofpacket,   --          .endofpacket
			src5_ready         => cmd_xbar_demux_001_src5_ready,         --      src5.ready
			src5_valid         => cmd_xbar_demux_001_src5_valid,         --          .valid
			src5_data          => cmd_xbar_demux_001_src5_data,          --          .data
			src5_channel       => cmd_xbar_demux_001_src5_channel,       --          .channel
			src5_startofpacket => cmd_xbar_demux_001_src5_startofpacket, --          .startofpacket
			src5_endofpacket   => cmd_xbar_demux_001_src5_endofpacket,   --          .endofpacket
			src6_ready         => cmd_xbar_demux_001_src6_ready,         --      src6.ready
			src6_valid         => cmd_xbar_demux_001_src6_valid,         --          .valid
			src6_data          => cmd_xbar_demux_001_src6_data,          --          .data
			src6_channel       => cmd_xbar_demux_001_src6_channel,       --          .channel
			src6_startofpacket => cmd_xbar_demux_001_src6_startofpacket, --          .startofpacket
			src6_endofpacket   => cmd_xbar_demux_001_src6_endofpacket,   --          .endofpacket
			src7_ready         => cmd_xbar_demux_001_src7_ready,         --      src7.ready
			src7_valid         => cmd_xbar_demux_001_src7_valid,         --          .valid
			src7_data          => cmd_xbar_demux_001_src7_data,          --          .data
			src7_channel       => cmd_xbar_demux_001_src7_channel,       --          .channel
			src7_startofpacket => cmd_xbar_demux_001_src7_startofpacket, --          .startofpacket
			src7_endofpacket   => cmd_xbar_demux_001_src7_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux : component nios_system_cmd_xbar_mux
		port map (
			clk                 => external_clocks_sys_clk_clk,           --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_src_ready,                --       src.ready
			src_valid           => cmd_xbar_mux_src_valid,                --          .valid
			src_data            => cmd_xbar_mux_src_data,                 --          .data
			src_channel         => cmd_xbar_mux_src_channel,              --          .channel
			src_startofpacket   => cmd_xbar_mux_src_startofpacket,        --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_src_endofpacket,          --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src0_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src0_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src0_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src0_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src0_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src0_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src0_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src0_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src0_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src0_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src0_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src0_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_001 : component nios_system_cmd_xbar_mux
		port map (
			clk                 => external_clocks_sys_clk_clk,           --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_001_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_001_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_001_src_data,             --          .data
			src_channel         => cmd_xbar_mux_001_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_001_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_001_src_endofpacket,      --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src1_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src1_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src1_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src1_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src1_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src1_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src1_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src1_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src1_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src1_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src1_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux : component nios_system_rsp_xbar_demux
		port map (
			clk                => external_clocks_sys_clk_clk,       --       clk.clk
			reset              => rst_controller_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_src_ready,               --      sink.ready
			sink_channel       => id_router_src_channel,             --          .channel
			sink_data          => id_router_src_data,                --          .data
			sink_startofpacket => id_router_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_001 : component nios_system_rsp_xbar_demux
		port map (
			clk                => external_clocks_sys_clk_clk,           --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => width_adapter_001_src_ready,           --      sink.ready
			sink_channel       => width_adapter_001_src_channel,         --          .channel
			sink_data          => width_adapter_001_src_data,            --          .data
			sink_startofpacket => width_adapter_001_src_startofpacket,   --          .startofpacket
			sink_endofpacket   => width_adapter_001_src_endofpacket,     --          .endofpacket
			sink_valid(0)      => width_adapter_001_src_valid,           --          .valid
			src0_ready         => rsp_xbar_demux_001_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_001_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_001_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_001_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_001_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_001_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_001_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_001_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_001_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_001_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_001_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_001_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_002 : component nios_system_rsp_xbar_demux_002
		port map (
			clk                => external_clocks_sys_clk_clk,           --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_002_src_ready,               --      sink.ready
			sink_channel       => id_router_002_src_channel,             --          .channel
			sink_data          => id_router_002_src_data,                --          .data
			sink_startofpacket => id_router_002_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_002_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_002_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_002_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_002_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_002_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_002_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_002_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_002_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_003 : component nios_system_rsp_xbar_demux_002
		port map (
			clk                => external_clocks_sys_clk_clk,           --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_003_src_ready,               --      sink.ready
			sink_channel       => id_router_003_src_channel,             --          .channel
			sink_data          => id_router_003_src_data,                --          .data
			sink_startofpacket => id_router_003_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_003_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_003_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_003_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_003_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_003_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_003_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_003_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_003_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_004 : component nios_system_rsp_xbar_demux_002
		port map (
			clk                => external_clocks_sys_clk_clk,           --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_004_src_ready,               --      sink.ready
			sink_channel       => id_router_004_src_channel,             --          .channel
			sink_data          => id_router_004_src_data,                --          .data
			sink_startofpacket => id_router_004_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_004_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_004_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_004_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_004_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_004_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_004_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_004_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_004_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_005 : component nios_system_rsp_xbar_demux_002
		port map (
			clk                => external_clocks_sys_clk_clk,           --       clk.clk
			reset              => cpu_jtag_debug_module_reset_reset,     -- clk_reset.reset
			sink_ready         => id_router_005_src_ready,               --      sink.ready
			sink_channel       => id_router_005_src_channel,             --          .channel
			sink_data          => id_router_005_src_data,                --          .data
			sink_startofpacket => id_router_005_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_005_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_005_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_005_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_005_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_005_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_005_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_005_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_005_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_006 : component nios_system_rsp_xbar_demux_002
		port map (
			clk                => external_clocks_sys_clk_clk,           --       clk.clk
			reset              => cpu_jtag_debug_module_reset_reset,     -- clk_reset.reset
			sink_ready         => id_router_006_src_ready,               --      sink.ready
			sink_channel       => id_router_006_src_channel,             --          .channel
			sink_data          => id_router_006_src_data,                --          .data
			sink_startofpacket => id_router_006_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_006_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_006_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_006_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_006_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_006_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_006_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_006_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_006_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_007 : component nios_system_rsp_xbar_demux_002
		port map (
			clk                => external_clocks_sys_clk_clk,           --       clk.clk
			reset              => cpu_jtag_debug_module_reset_reset,     -- clk_reset.reset
			sink_ready         => id_router_007_src_ready,               --      sink.ready
			sink_channel       => id_router_007_src_channel,             --          .channel
			sink_data          => id_router_007_src_data,                --          .data
			sink_startofpacket => id_router_007_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_007_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_007_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_007_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_007_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_007_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_007_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_007_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_007_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_mux : component nios_system_rsp_xbar_mux
		port map (
			clk                 => external_clocks_sys_clk_clk,           --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => rsp_xbar_mux_src_ready,                --       src.ready
			src_valid           => rsp_xbar_mux_src_valid,                --          .valid
			src_data            => rsp_xbar_mux_src_data,                 --          .data
			src_channel         => rsp_xbar_mux_src_channel,              --          .channel
			src_startofpacket   => rsp_xbar_mux_src_startofpacket,        --          .startofpacket
			src_endofpacket     => rsp_xbar_mux_src_endofpacket,          --          .endofpacket
			sink0_ready         => rsp_xbar_demux_src0_ready,             --     sink0.ready
			sink0_valid         => rsp_xbar_demux_src0_valid,             --          .valid
			sink0_channel       => rsp_xbar_demux_src0_channel,           --          .channel
			sink0_data          => rsp_xbar_demux_src0_data,              --          .data
			sink0_startofpacket => rsp_xbar_demux_src0_startofpacket,     --          .startofpacket
			sink0_endofpacket   => rsp_xbar_demux_src0_endofpacket,       --          .endofpacket
			sink1_ready         => rsp_xbar_demux_001_src0_ready,         --     sink1.ready
			sink1_valid         => rsp_xbar_demux_001_src0_valid,         --          .valid
			sink1_channel       => rsp_xbar_demux_001_src0_channel,       --          .channel
			sink1_data          => rsp_xbar_demux_001_src0_data,          --          .data
			sink1_startofpacket => rsp_xbar_demux_001_src0_startofpacket, --          .startofpacket
			sink1_endofpacket   => rsp_xbar_demux_001_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_mux_001 : component nios_system_rsp_xbar_mux_001
		port map (
			clk                 => external_clocks_sys_clk_clk,           --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => rsp_xbar_mux_001_src_ready,            --       src.ready
			src_valid           => rsp_xbar_mux_001_src_valid,            --          .valid
			src_data            => rsp_xbar_mux_001_src_data,             --          .data
			src_channel         => rsp_xbar_mux_001_src_channel,          --          .channel
			src_startofpacket   => rsp_xbar_mux_001_src_startofpacket,    --          .startofpacket
			src_endofpacket     => rsp_xbar_mux_001_src_endofpacket,      --          .endofpacket
			sink0_ready         => rsp_xbar_demux_src1_ready,             --     sink0.ready
			sink0_valid         => rsp_xbar_demux_src1_valid,             --          .valid
			sink0_channel       => rsp_xbar_demux_src1_channel,           --          .channel
			sink0_data          => rsp_xbar_demux_src1_data,              --          .data
			sink0_startofpacket => rsp_xbar_demux_src1_startofpacket,     --          .startofpacket
			sink0_endofpacket   => rsp_xbar_demux_src1_endofpacket,       --          .endofpacket
			sink1_ready         => rsp_xbar_demux_001_src1_ready,         --     sink1.ready
			sink1_valid         => rsp_xbar_demux_001_src1_valid,         --          .valid
			sink1_channel       => rsp_xbar_demux_001_src1_channel,       --          .channel
			sink1_data          => rsp_xbar_demux_001_src1_data,          --          .data
			sink1_startofpacket => rsp_xbar_demux_001_src1_startofpacket, --          .startofpacket
			sink1_endofpacket   => rsp_xbar_demux_001_src1_endofpacket,   --          .endofpacket
			sink2_ready         => rsp_xbar_demux_002_src0_ready,         --     sink2.ready
			sink2_valid         => rsp_xbar_demux_002_src0_valid,         --          .valid
			sink2_channel       => rsp_xbar_demux_002_src0_channel,       --          .channel
			sink2_data          => rsp_xbar_demux_002_src0_data,          --          .data
			sink2_startofpacket => rsp_xbar_demux_002_src0_startofpacket, --          .startofpacket
			sink2_endofpacket   => rsp_xbar_demux_002_src0_endofpacket,   --          .endofpacket
			sink3_ready         => rsp_xbar_demux_003_src0_ready,         --     sink3.ready
			sink3_valid         => rsp_xbar_demux_003_src0_valid,         --          .valid
			sink3_channel       => rsp_xbar_demux_003_src0_channel,       --          .channel
			sink3_data          => rsp_xbar_demux_003_src0_data,          --          .data
			sink3_startofpacket => rsp_xbar_demux_003_src0_startofpacket, --          .startofpacket
			sink3_endofpacket   => rsp_xbar_demux_003_src0_endofpacket,   --          .endofpacket
			sink4_ready         => rsp_xbar_demux_004_src0_ready,         --     sink4.ready
			sink4_valid         => rsp_xbar_demux_004_src0_valid,         --          .valid
			sink4_channel       => rsp_xbar_demux_004_src0_channel,       --          .channel
			sink4_data          => rsp_xbar_demux_004_src0_data,          --          .data
			sink4_startofpacket => rsp_xbar_demux_004_src0_startofpacket, --          .startofpacket
			sink4_endofpacket   => rsp_xbar_demux_004_src0_endofpacket,   --          .endofpacket
			sink5_ready         => rsp_xbar_demux_005_src0_ready,         --     sink5.ready
			sink5_valid         => rsp_xbar_demux_005_src0_valid,         --          .valid
			sink5_channel       => rsp_xbar_demux_005_src0_channel,       --          .channel
			sink5_data          => rsp_xbar_demux_005_src0_data,          --          .data
			sink5_startofpacket => rsp_xbar_demux_005_src0_startofpacket, --          .startofpacket
			sink5_endofpacket   => rsp_xbar_demux_005_src0_endofpacket,   --          .endofpacket
			sink6_ready         => rsp_xbar_demux_006_src0_ready,         --     sink6.ready
			sink6_valid         => rsp_xbar_demux_006_src0_valid,         --          .valid
			sink6_channel       => rsp_xbar_demux_006_src0_channel,       --          .channel
			sink6_data          => rsp_xbar_demux_006_src0_data,          --          .data
			sink6_startofpacket => rsp_xbar_demux_006_src0_startofpacket, --          .startofpacket
			sink6_endofpacket   => rsp_xbar_demux_006_src0_endofpacket,   --          .endofpacket
			sink7_ready         => rsp_xbar_demux_007_src0_ready,         --     sink7.ready
			sink7_valid         => rsp_xbar_demux_007_src0_valid,         --          .valid
			sink7_channel       => rsp_xbar_demux_007_src0_channel,       --          .channel
			sink7_data          => rsp_xbar_demux_007_src0_data,          --          .data
			sink7_startofpacket => rsp_xbar_demux_007_src0_startofpacket, --          .startofpacket
			sink7_endofpacket   => rsp_xbar_demux_007_src0_endofpacket    --          .endofpacket
		);

	width_adapter : component nios_system_width_adapter
		generic map (
			IN_PKT_ADDR_H                 => 64,
			IN_PKT_ADDR_L                 => 36,
			IN_PKT_DATA_H                 => 31,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 35,
			IN_PKT_BYTEEN_L               => 32,
			IN_PKT_BYTE_CNT_H             => 73,
			IN_PKT_BYTE_CNT_L             => 71,
			IN_PKT_TRANS_COMPRESSED_READ  => 65,
			IN_PKT_BURSTWRAP_H            => 76,
			IN_PKT_BURSTWRAP_L            => 74,
			IN_PKT_BURST_SIZE_H           => 79,
			IN_PKT_BURST_SIZE_L           => 77,
			IN_PKT_RESPONSE_STATUS_H      => 101,
			IN_PKT_RESPONSE_STATUS_L      => 100,
			IN_PKT_TRANS_EXCLUSIVE        => 70,
			IN_PKT_BURST_TYPE_H           => 81,
			IN_PKT_BURST_TYPE_L           => 80,
			IN_ST_DATA_W                  => 102,
			OUT_PKT_ADDR_H                => 46,
			OUT_PKT_ADDR_L                => 18,
			OUT_PKT_DATA_H                => 15,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 17,
			OUT_PKT_BYTEEN_L              => 16,
			OUT_PKT_BYTE_CNT_H            => 55,
			OUT_PKT_BYTE_CNT_L            => 53,
			OUT_PKT_TRANS_COMPRESSED_READ => 47,
			OUT_PKT_BURST_SIZE_H          => 61,
			OUT_PKT_BURST_SIZE_L          => 59,
			OUT_PKT_RESPONSE_STATUS_H     => 83,
			OUT_PKT_RESPONSE_STATUS_L     => 82,
			OUT_PKT_TRANS_EXCLUSIVE       => 52,
			OUT_PKT_BURST_TYPE_H          => 63,
			OUT_PKT_BURST_TYPE_L          => 62,
			OUT_ST_DATA_W                 => 84,
			ST_CHANNEL_W                  => 8,
			OPTIMIZE_FOR_RSP              => 0,
			RESPONSE_PATH                 => 0
		)
		port map (
			clk                  => external_clocks_sys_clk_clk,        --       clk.clk
			reset                => rst_controller_reset_out_reset,     -- clk_reset.reset
			in_valid             => cmd_xbar_mux_001_src_valid,         --      sink.valid
			in_channel           => cmd_xbar_mux_001_src_channel,       --          .channel
			in_startofpacket     => cmd_xbar_mux_001_src_startofpacket, --          .startofpacket
			in_endofpacket       => cmd_xbar_mux_001_src_endofpacket,   --          .endofpacket
			in_ready             => cmd_xbar_mux_001_src_ready,         --          .ready
			in_data              => cmd_xbar_mux_001_src_data,          --          .data
			out_endofpacket      => width_adapter_src_endofpacket,      --       src.endofpacket
			out_data             => width_adapter_src_data,             --          .data
			out_channel          => width_adapter_src_channel,          --          .channel
			out_valid            => width_adapter_src_valid,            --          .valid
			out_ready            => width_adapter_src_ready,            --          .ready
			out_startofpacket    => width_adapter_src_startofpacket,    --          .startofpacket
			in_command_size_data => "000"                               -- (terminated)
		);

	width_adapter_001 : component nios_system_width_adapter_001
		generic map (
			IN_PKT_ADDR_H                 => 46,
			IN_PKT_ADDR_L                 => 18,
			IN_PKT_DATA_H                 => 15,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 17,
			IN_PKT_BYTEEN_L               => 16,
			IN_PKT_BYTE_CNT_H             => 55,
			IN_PKT_BYTE_CNT_L             => 53,
			IN_PKT_TRANS_COMPRESSED_READ  => 47,
			IN_PKT_BURSTWRAP_H            => 58,
			IN_PKT_BURSTWRAP_L            => 56,
			IN_PKT_BURST_SIZE_H           => 61,
			IN_PKT_BURST_SIZE_L           => 59,
			IN_PKT_RESPONSE_STATUS_H      => 83,
			IN_PKT_RESPONSE_STATUS_L      => 82,
			IN_PKT_TRANS_EXCLUSIVE        => 52,
			IN_PKT_BURST_TYPE_H           => 63,
			IN_PKT_BURST_TYPE_L           => 62,
			IN_ST_DATA_W                  => 84,
			OUT_PKT_ADDR_H                => 64,
			OUT_PKT_ADDR_L                => 36,
			OUT_PKT_DATA_H                => 31,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 35,
			OUT_PKT_BYTEEN_L              => 32,
			OUT_PKT_BYTE_CNT_H            => 73,
			OUT_PKT_BYTE_CNT_L            => 71,
			OUT_PKT_TRANS_COMPRESSED_READ => 65,
			OUT_PKT_BURST_SIZE_H          => 79,
			OUT_PKT_BURST_SIZE_L          => 77,
			OUT_PKT_RESPONSE_STATUS_H     => 101,
			OUT_PKT_RESPONSE_STATUS_L     => 100,
			OUT_PKT_TRANS_EXCLUSIVE       => 70,
			OUT_PKT_BURST_TYPE_H          => 81,
			OUT_PKT_BURST_TYPE_L          => 80,
			OUT_ST_DATA_W                 => 102,
			ST_CHANNEL_W                  => 8,
			OPTIMIZE_FOR_RSP              => 1,
			RESPONSE_PATH                 => 1
		)
		port map (
			clk                  => external_clocks_sys_clk_clk,         --       clk.clk
			reset                => rst_controller_reset_out_reset,      -- clk_reset.reset
			in_valid             => id_router_001_src_valid,             --      sink.valid
			in_channel           => id_router_001_src_channel,           --          .channel
			in_startofpacket     => id_router_001_src_startofpacket,     --          .startofpacket
			in_endofpacket       => id_router_001_src_endofpacket,       --          .endofpacket
			in_ready             => id_router_001_src_ready,             --          .ready
			in_data              => id_router_001_src_data,              --          .data
			out_endofpacket      => width_adapter_001_src_endofpacket,   --       src.endofpacket
			out_data             => width_adapter_001_src_data,          --          .data
			out_channel          => width_adapter_001_src_channel,       --          .channel
			out_valid            => width_adapter_001_src_valid,         --          .valid
			out_ready            => width_adapter_001_src_ready,         --          .ready
			out_startofpacket    => width_adapter_001_src_startofpacket, --          .startofpacket
			in_command_size_data => "000"                                -- (terminated)
		);

	irq_mapper : component nios_system_irq_mapper
		port map (
			clk           => external_clocks_sys_clk_clk,    --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			sender_irq    => cpu_d_irq_irq                   --    sender.irq
		);

	reset_n_ports_inv <= not reset_n;

	sdram_s1_translator_avalon_anti_slave_0_write_ports_inv <= not sdram_s1_translator_avalon_anti_slave_0_write;

	sdram_s1_translator_avalon_anti_slave_0_read_ports_inv <= not sdram_s1_translator_avalon_anti_slave_0_read;

	sdram_s1_translator_avalon_anti_slave_0_byteenable_ports_inv <= not sdram_s1_translator_avalon_anti_slave_0_byteenable;

	interval_timer_s1_translator_avalon_anti_slave_0_write_ports_inv <= not interval_timer_s1_translator_avalon_anti_slave_0_write;

	jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write_ports_inv <= not jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write;

	jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read_ports_inv <= not jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of nios_system
